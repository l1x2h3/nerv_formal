`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [31:0] PI_io_tlb_Anotherread_2_data;
  reg [31:0] PI_io_tlb_Anotherread_0_data;
  reg [31:0] PI_io_inst;
  wire [0:0] PI_clock = clock;
  reg [31:0] PI_irq;
  reg [0:0] PI_stall;
  reg [31:0] PI_io_tlb_Anotherread_1_data;
  reg [0:0] PI_reset;
  reg [31:0] PI_io_mem_read_data;
  reg [0:0] PI_io_valid;
  top_formal UUT (
    .io_tlb_Anotherread_2_data(PI_io_tlb_Anotherread_2_data),
    .io_tlb_Anotherread_0_data(PI_io_tlb_Anotherread_0_data),
    .io_inst(PI_io_inst),
    .clock(PI_clock),
    .irq(PI_irq),
    .stall(PI_stall),
    .io_tlb_Anotherread_1_data(PI_io_tlb_Anotherread_1_data),
    .reset(PI_reset),
    .io_mem_read_data(PI_io_mem_read_data),
    .io_valid(PI_io_valid)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18570  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18600  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18882  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18900  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18912  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18918  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$18924  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18574  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18580  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18586  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18592  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18598  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18604  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18610  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18616  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18622  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18628  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18634  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18640  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18646  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18652  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18658  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18664  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18670  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18676  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18682  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18688  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18694  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18700  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18706  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18712  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18718  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18724  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18730  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18736  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18742  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18748  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18754  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18760  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18766  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18772  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18778  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18784  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18790  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18796  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18802  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18808  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18814  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18820  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18826  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18832  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18838  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18844  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18850  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18856  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18862  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18868  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18874  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18880  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18886  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18892  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18898  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18904  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18910  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18916  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18922  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$18928  = 1'b1;
    UUT.checker_inst.checker_.LoadQueue.queue_q.deq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.LoadQueue.queue_q.enq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.LoadQueue.queue_q.maybe_full = 1'b0;
    UUT.checker_inst.checker_.StoreQueue.queue_q.deq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.StoreQueue.queue_q.enq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.StoreQueue.queue_q.maybe_full = 1'b0;
    UUT.checker_inst.checker_.TLBLoadQueue_0.queue_q.deq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.TLBLoadQueue_0.queue_q.enq_ptr_value = 1'b1;
    UUT.checker_inst.checker_.TLBLoadQueue_0.queue_q.maybe_full = 1'b0;
    UUT.checker_inst.checker_.TLBLoadQueue_1.queue_q.deq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.TLBLoadQueue_1.queue_q.enq_ptr_value = 1'b1;
    UUT.checker_inst.checker_.TLBLoadQueue_1.queue_q.maybe_full = 1'b0;
    UUT.checker_inst.checker_.TLBLoadQueue_2.queue_q.deq_ptr_value = 1'b0;
    UUT.checker_inst.checker_.TLBLoadQueue_2.queue_q.enq_ptr_value = 1'b1;
    UUT.checker_inst.checker_.TLBLoadQueue_2.queue_q.maybe_full = 1'b0;
    UUT.checker_inst.checker_.specCore.state_csr_IALIGN = 8'b00000000;
    UUT.checker_inst.checker_.specCore.state_csr_MXLEN = 8'b00000000;
    UUT.checker_inst.checker_.specCore.state_csr_marchid = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mcause = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mcounteren = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_medeleg = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mepc = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mhartid = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mie = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mimpid = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mip = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_misa = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mscratch = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mstatus = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mtval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mtvec = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mvendorid = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_satp = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_scause = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_sepc = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_stvec = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_internal_privilegeMode = 2'b00;
    UUT.checker_inst.checker_.specCore.state_pc = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_10 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_12 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_13 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_14 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_15 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_16 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_17 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_18 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_19 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_2 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_20 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_21 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_22 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_24 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_25 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_26 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_27 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_28 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_29 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_3 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_30 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_31 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_4 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_5 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_6 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_7 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_8 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_9 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.csr_marchid = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mcause = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mcounteren = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mepc = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mhartid = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mie = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mimpid = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mip = 32'b00000000000000000000000000000000;
    UUT.dut.csr_misa = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mscratch = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mstatus = 32'b00000000000000000001100000000000;
    UUT.dut.csr_mtval = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mtvec = 32'b00000000000000000000000000000000;
    UUT.dut.csr_mvendorid = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_custom_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_hpm_counter_value = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_hpm_counterh_value = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_hpm_event_value = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mcause_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mepc_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mie_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mip_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_misa_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mscratch_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mstatus_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mstatush_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mtval_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.csr_mtvec_value = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.mem_rd_enable_q = 1'b0;
    UUT.dut.nerv_inst.mem_rd_func_q = 5'b00000;
    UUT.dut.nerv_inst.mem_rd_reg_q = 5'b10000;
    UUT.dut.nerv_inst.mem_wr_enable_q = 1'b0;
    UUT.dut.nerv_inst.next_rvfi_intr = 1'b0;
    UUT.dut.nerv_inst.pc = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.reset_q = 1'b0;
    UUT.dut.nerv_inst.rvfi_csr_custom_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_ro_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_ro_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_ro_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_ro_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_custom_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_marchid_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_marchid_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_marchid_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_marchid_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcause_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcause_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcause_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcause_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mconfigptr_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mconfigptr_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mconfigptr_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mconfigptr_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycle_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycle_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycle_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycle_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycleh_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycleh_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycleh_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mcycleh_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mepc_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mepc_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mepc_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mepc_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhartid_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhartid_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhartid_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhartid_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter10h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter11h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter12h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter13h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter14h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter15h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter16h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter17h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter18h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter19h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter20h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter21h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter22h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter23h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter24h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter25h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter26h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter27h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter28h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter29h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter30h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter31h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter3h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter4h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter5h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter6h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter7h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter8h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9h_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9h_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9h_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmcounter9h_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent10_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent10_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent10_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent10_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent11_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent11_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent11_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent11_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent12_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent12_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent12_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent12_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent13_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent13_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent13_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent13_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent14_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent14_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent14_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent14_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent15_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent15_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent15_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent15_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent16_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent16_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent16_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent16_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent17_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent17_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent17_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent17_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent18_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent18_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent18_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent18_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent19_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent19_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent19_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent19_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent20_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent20_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent20_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent20_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent21_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent21_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent21_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent21_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent22_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent22_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent22_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent22_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent23_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent23_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent23_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent23_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent24_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent24_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent24_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent24_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent25_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent25_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent25_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent25_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent26_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent26_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent26_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent26_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent27_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent27_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent27_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent27_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent28_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent28_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent28_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent28_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent29_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent29_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent29_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent29_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent30_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent30_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent30_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent30_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent31_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent31_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent31_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent31_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent3_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent3_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent3_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent3_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent4_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent4_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent4_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent4_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent5_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent5_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent5_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent5_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent6_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent6_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent6_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent6_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent7_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent7_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent7_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent7_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent8_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent8_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent8_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent8_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent9_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent9_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent9_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mhpmevent9_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mie_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mie_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mie_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mie_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mimpid_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mimpid_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mimpid_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mimpid_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstret_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstret_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstret_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstret_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstreth_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstreth_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstreth_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_minstreth_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mip_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mip_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mip_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mip_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_misa_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_misa_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_misa_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_misa_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mscratch_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mscratch_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mscratch_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mscratch_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatus_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatus_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatus_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatus_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatush_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatush_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatush_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mstatush_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtval_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtval_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtval_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtval_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtvec_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtvec_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtvec_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mtvec_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mvendorid_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mvendorid_rmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mvendorid_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_csr_mvendorid_wmask = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_halt = 1'b0;
    UUT.dut.nerv_inst.rvfi_insn = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_intr = 1'b0;
    UUT.dut.nerv_inst.rvfi_ixl = 2'b00;
    UUT.dut.nerv_inst.rvfi_mem_addr = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_mem_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_mem_rmask = 4'b0000;
    UUT.dut.nerv_inst.rvfi_mem_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_mem_wmask = 4'b0000;
    UUT.dut.nerv_inst.rvfi_mode = 2'b00;
    UUT.dut.nerv_inst.rvfi_order = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_pc_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_pc_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_rd_addr = 5'b00000;
    UUT.dut.nerv_inst.rvfi_rd_wdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_rs1_addr = 5'b00000;
    UUT.dut.nerv_inst.rvfi_rs1_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_rs2_addr = 5'b00000;
    UUT.dut.nerv_inst.rvfi_rs2_rdata = 32'b00000000000000000000000000000000;
    UUT.dut.nerv_inst.rvfi_trap = 1'b0;
    UUT.dut.nerv_inst.rvfi_valid = 1'b0;
    UUT.checker_inst.checker_.LoadQueue.queue_q.ram_addr[1'b0] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.LoadQueue.queue_q.ram_data[1'b0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.LoadQueue.queue_q.ram_memWidth[1'b0] = 7'b1000000;
    UUT.checker_inst.checker_.StoreQueue.queue_q.ram_addr[1'b0] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.StoreQueue.queue_q.ram_data[1'b0] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.StoreQueue.queue_q.ram_memWidth[1'b0] = 7'b1000000;
    UUT.checker_inst.checker_.TLBLoadQueue_0.queue_q.ram_addr[1'b0] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.TLBLoadQueue_0.queue_q.ram_data[1'b0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.TLBLoadQueue_1.queue_q.ram_addr[1'b0] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.TLBLoadQueue_1.queue_q.ram_data[1'b0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.TLBLoadQueue_2.queue_q.ram_addr[1'b0] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.checker_inst.checker_.TLBLoadQueue_2.queue_q.ram_data[1'b0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.nerv_inst.regfile[5'b00000] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11111] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11110] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11101] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11100] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11011] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11010] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11001] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b11000] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10111] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10110] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10101] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10100] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10011] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10010] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10001] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b10000] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01111] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01110] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01101] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01100] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01011] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01010] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01001] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b01000] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00111] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00110] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00101] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00100] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00011] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00010] = 32'b00000000000000000000000000000000;
    UUT.dut.regfile[5'b00001] = 32'b00000000000000000000000000000000;

    // state 0
    PI_io_tlb_Anotherread_2_data = 32'b00000000000000000000000000000000;
    PI_io_tlb_Anotherread_0_data = 32'b00000000000000000000000000000000;
    PI_io_inst = 32'b00000000000000000000000000000000;
    PI_irq = 32'b00000000000000000000000000000000;
    PI_stall = 1'b0;
    PI_io_tlb_Anotherread_1_data = 32'b00000000000000000000000000000000;
    PI_reset = 1'b0;
    PI_io_mem_read_data = 32'b00000000000000000000000000000000;
    PI_io_valid = 1'b0;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_io_tlb_Anotherread_2_data <= 32'b00000000000000000000000000000000;
      PI_io_tlb_Anotherread_0_data <= 32'b00000000000000000000000000000000;
      PI_io_inst <= 32'b00000000000000000000000000000000;
      PI_irq <= 32'b00000000000000000000000000000000;
      PI_stall <= 1'b0;
      PI_io_tlb_Anotherread_1_data <= 32'b00000000000000000000000000000000;
      PI_reset <= 1'b0;
      PI_io_mem_read_data <= 32'b00000000000000000000000000000000;
      PI_io_valid <= 1'b0;
    end

    genclock <= cycle < 1;
    cycle <= cycle + 1;
  end
endmodule
