module RiscvTrans(
  input         clock,
  input         reset,
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_iFetchpc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [1:0]  io_now_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [1:0]  io_next_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
);
  wire  _exceptionVec_WIRE_5 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_5 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_7 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_7 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_1 = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_13 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_13 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_2 = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_15 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_15 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_3 = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] inst = io_valid ? io_inst : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_6103 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _T_426 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_427 = 32'h5003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_444 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _T_1081 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1082 = 32'h7073 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_1083 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_65 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_1040 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1041 = 32'h6073 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_1042 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_64 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_1006 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1007 = 32'h5073 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_1008 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_63 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_966 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_967 = 32'h3073 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_968 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_62 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_926 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_927 = 32'h2073 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_928 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_61 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_893 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_894 = 32'h1073 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_895 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_60 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_887 = inst & 32'hfe007fff; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_888 = 32'h12000073 == _T_887; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_889 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_59 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_881 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_882 = 32'h10500073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_883 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_58 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_874 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_875 = 32'h30200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_876 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_57 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_867 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_868 = 32'h10200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_869 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_56 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_860 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_861 = 32'h2007033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_862 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_863 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_55 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_853 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_854 = 32'h2006033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_855 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_856 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_54 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_846 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_847 = 32'h2005033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_848 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_849 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_53 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_839 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_840 = 32'h2004033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_841 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_842 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_52 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_832 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_833 = 32'h2003033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_834 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_835 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_51 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_825 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_826 = 32'h2002033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_827 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_828 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_50 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_818 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_819 = 32'h2001033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_820 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_821 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_49 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_811 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_812 = 32'h2000033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_813 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_814 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_48 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_804 = inst & 32'hef83; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_805 = 32'h1 == _T_804; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [15:0] _T_806 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_807 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_808 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_47 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_760 = inst & 32'hf003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_761 = 32'h9002 == _T_760; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_762 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_763 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire [4:0] _T_764 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 76:112]
  wire  _T_765 = inst[6:2] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 76:119]
  wire  _T_766 = _T_763 & inst[6:2] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 76:105]
  wire  _T_767 = 32'h9002 == _T_760 & _T_766; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_768 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:97]
  wire [11:0] _T_769 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_46 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_748 = inst & 32'hf003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_749 = 32'h8002 == _T_760; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_750 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_751 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire [4:0] _T_752 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 73:112]
  wire  _T_753 = inst[6:2] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 73:119]
  wire  _T_754 = _T_763 & _T_765; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 73:105]
  wire  _T_755 = 32'h8002 == _T_760 & _T_766; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_756 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:97]
  wire [11:0] _T_757 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_45 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_690 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_691 = 32'h2 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_692 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_693 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_694 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 15:22]
  wire  _T_695 = ~inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 15:27]
  wire  _T_696 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:19]
  wire [4:0] _T_697 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:29]
  wire [5:0] _T_698 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:14]
  wire  _T_699 = _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:37]
  wire  _T_700 = _T_695 & _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:8]
  wire  _T_701 = _T_763 & _T_700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 65:105]
  wire  _T_702 = 32'h2 == _T_690 & _T_701; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_703 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_704 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_705 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_44 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_668 = inst & 32'hef83; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_669 = 32'h6101 == _T_804; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_670 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:59]
  wire [4:0] _T_671 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:69]
  wire [5:0] _T_672 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:54]
  wire  _T_673 = _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:77]
  wire  _T_674 = 32'h6101 == _T_804 & _T_699; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_675 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_676 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_677 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_43 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_653 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_654 = 32'h1 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_655 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_656 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_657 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:59]
  wire [4:0] _T_658 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:69]
  wire [5:0] _T_659 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:54]
  wire  _T_660 = _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:77]
  wire  _T_661 = _T_763 & _T_699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 39:107]
  wire  _T_662 = 32'h1 == _T_690 & _T_661; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_663 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_664 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_665 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_42 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_635 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_636 = 32'h6001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_637 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_638 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire [4:0] _T_639 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 44:114]
  wire  _T_640 = inst[11:7] != 5'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 44:122]
  wire  _T_641 = _T_763 & inst[11:7] != 5'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 44:107]
  wire  _T_642 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:59]
  wire [4:0] _T_643 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:69]
  wire [5:0] _T_644 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:54]
  wire  _T_645 = _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 12:77]
  wire  _T_646 = _T_763 & inst[11:7] != 5'h2 & _T_699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 44:130]
  wire  _T_647 = 32'h6001 == _T_690 & _T_646; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_648 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_649 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_650 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_41 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_625 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_626 = 32'h4001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_627 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_628 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_629 = 32'h4001 == _T_690 & _T_763; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_630 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_631 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_632 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_40 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_598 = inst & 32'hf07f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_599 = 32'h9002 == _T_598; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_600 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_601 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_602 = 32'h9002 == _T_598 & _T_763; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_603 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:97]
  wire [11:0] _T_604 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_39 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_589 = inst & 32'hf07f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_590 = 32'h8002 == _T_598; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_591 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_592 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_593 = 32'h8002 == _T_598 & _T_763; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_594 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:97]
  wire [11:0] _T_595 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_38 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_538 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_539 = 32'h4002 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [4:0] _T_540 = inst[11:7]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:55]
  wire  _T_541 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_542 = 32'h4002 == _T_690 & _T_763; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [15:0] _T_543 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:97]
  wire [12:0] _T_544 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_545 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_37 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_532 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_533 = 32'hf == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_534 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_36 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_523 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_524 = 32'h73 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_525 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_35 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_517 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_518 = 32'h100073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_519 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_34 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_493 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_494 = 32'h2023 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_495 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_496 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_33 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_469 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_470 = 32'h1023 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_471 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_472 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_32 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_446 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_447 = 32'h23 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_448 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_449 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_31 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [19:0] _T_428 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_30 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_407 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_408 = 32'h4003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_409 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_29 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_387 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_388 = 32'h2003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_389 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_28 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_367 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_368 = 32'h1003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_369 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_27 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_347 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_348 = 32'h3 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_349 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_26 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_320 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_321 = 32'h7063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_322 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_323 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_324 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_25 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_291 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_292 = 32'h5063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_293 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_294 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_295 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_24 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_264 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_265 = 32'h6063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_266 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_267 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_268 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_23 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_235 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_236 = 32'h4063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_237 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_238 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_239 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_22 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_208 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_209 = 32'h1063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_210 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_211 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_212 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_21 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_181 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_182 = 32'h63 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_183 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_184 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_185 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_20 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_156 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_157 = 32'h67 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_158 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_19 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_125 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_126 = 32'h40005033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_127 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_128 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_18 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_118 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_119 = 32'h40000033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_120 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_121 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_17 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_111 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_112 = 32'h5033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_113 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_114 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_16 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_104 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_105 = 32'h1033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_106 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_107 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_15 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_97 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_98 = 32'h4033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_99 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_100 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_14 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_90 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_91 = 32'h6033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_92 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_93 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_13 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_83 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_84 = 32'h7033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_85 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_86 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_12 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_76 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_77 = 32'h3033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_78 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_79 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_11 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_69 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_70 = 32'h2033 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_71 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_72 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_10 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_62 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_63 = 32'h33 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_64 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_65 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_9 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_48 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_49 = 32'h40005013 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [19:0] _T_50 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_8 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_42 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_43 = 32'h5013 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [19:0] _T_44 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_7 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_36 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_37 = 32'h1013 == _T_860; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [19:0] _T_38 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_6 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_30 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_31 = 32'h4013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_32 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_5 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_24 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_25 = 32'h6013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_26 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_4 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_18 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_19 = 32'h7013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_20 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_3 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_12 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_13 = 32'h3013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_14 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_2 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_6 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_7 = 32'h2013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_8 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_1 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1 = 32'h13 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_2 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_66 = _T_1 ? inst[19:15] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [4:0] _GEN_137 = _T_7 ? inst[19:15] : _GEN_66; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_208 = _T_13 ? inst[19:15] : _GEN_137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_279 = _T_19 ? inst[19:15] : _GEN_208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_350 = _T_25 ? inst[19:15] : _GEN_279; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_421 = _T_31 ? inst[19:15] : _GEN_350; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_492 = _T_37 ? inst[19:15] : _GEN_421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_563 = _T_43 ? inst[19:15] : _GEN_492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_634 = _T_49 ? inst[19:15] : _GEN_563; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_876 = _T_63 ? inst[19:15] : _GEN_634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_947 = _T_70 ? inst[19:15] : _GEN_876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1018 = _T_77 ? inst[19:15] : _GEN_947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1089 = _T_84 ? inst[19:15] : _GEN_1018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1160 = _T_91 ? inst[19:15] : _GEN_1089; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1231 = _T_98 ? inst[19:15] : _GEN_1160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1302 = _T_105 ? inst[19:15] : _GEN_1231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1373 = _T_112 ? inst[19:15] : _GEN_1302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1444 = _T_119 ? inst[19:15] : _GEN_1373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1515 = _T_126 ? inst[19:15] : _GEN_1444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1736 = _T_157 ? inst[19:15] : _GEN_1515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1792 = _T_182 ? inst[19:15] : _GEN_1736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1817 = _T_209 ? inst[19:15] : _GEN_1792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1842 = _T_236 ? inst[19:15] : _GEN_1817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1867 = _T_265 ? inst[19:15] : _GEN_1842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1892 = _T_292 ? inst[19:15] : _GEN_1867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1917 = _T_321 ? inst[19:15] : _GEN_1892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1999 = _T_348 ? inst[19:15] : _GEN_1917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2112 = _T_368 ? inst[19:15] : _GEN_1999; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2225 = _T_388 ? inst[19:15] : _GEN_2112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2303 = _T_408 ? inst[19:15] : _GEN_2225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2416 = _T_427 ? inst[19:15] : _GEN_2303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2463 = _T_447 ? inst[19:15] : _GEN_2416; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2483 = _T_470 ? inst[19:15] : _GEN_2463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2503 = _T_494 ? inst[19:15] : _GEN_2483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2516 = _T_518 ? inst[19:15] : _GEN_2503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2534 = _T_524 ? inst[19:15] : _GEN_2516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2545 = _T_533 ? inst[19:15] : _GEN_2534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2585 = _T_542 ? inst[11:7] : _GEN_2545; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2835 = _T_593 ? inst[11:7] : _GEN_2585; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2843 = _T_602 ? inst[11:7] : _GEN_2835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2973 = _T_629 ? inst[11:7] : _GEN_2843; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3045 = _T_647 ? inst[11:7] : _GEN_2973; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3148 = _T_662 ? inst[11:7] : _GEN_3045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3187 = _T_674 ? inst[11:7] : _GEN_3148; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3296 = _T_702 ? inst[11:7] : _GEN_3187; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3679 = _T_755 ? inst[11:7] : _GEN_3296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3749 = _T_767 ? inst[11:7] : _GEN_3679; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4328 = _T_805 ? inst[11:7] : _GEN_3749; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4367 = _T_812 ? inst[19:15] : _GEN_4328; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4438 = _T_819 ? inst[19:15] : _GEN_4367; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4509 = _T_826 ? inst[19:15] : _GEN_4438; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4580 = _T_833 ? inst[19:15] : _GEN_4509; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4651 = _T_840 ? inst[19:15] : _GEN_4580; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4722 = _T_847 ? inst[19:15] : _GEN_4651; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4793 = _T_854 ? inst[19:15] : _GEN_4722; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4864 = _T_861 ? inst[19:15] : _GEN_4793; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4913 = _T_868 ? inst[19:15] : _GEN_4864; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4934 = _T_875 ? inst[19:15] : _GEN_4913; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4948 = _T_882 ? inst[19:15] : _GEN_4934; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4955 = _T_888 ? inst[19:15] : _GEN_4948; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5098 = _T_894 ? inst[19:15] : _GEN_4955; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5270 = _T_927 ? inst[19:15] : _GEN_5098; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5442 = _T_967 ? inst[19:15] : _GEN_5270; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5630 = _T_1007 ? inst[19:15] : _GEN_5442; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5802 = _T_1041 ? inst[19:15] : _GEN_5630; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5974 = _T_1082 ? inst[19:15] : _GEN_5802; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs1 = io_valid ? _GEN_5974 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [4:0] _GEN_6106 = rs1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [31:0] now_reg_31 = io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_30 = io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_29 = io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_28 = io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_27 = io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_26 = io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_25 = io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_24 = io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_23 = io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_22 = io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_21 = io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_20 = io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_19 = io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_18 = io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_17 = io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_16 = io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_15 = io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_14 = io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_13 = io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_12 = io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_11 = io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_10 = io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_9 = io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_8 = io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_7 = io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_6 = io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_5 = io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_4 = io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_3 = io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_2 = io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_1 = io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_0 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_0 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_1 = 5'h1 == rs1 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_2 = 5'h2 == rs1 ? io_now_reg_2 : _GEN_1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_3 = 5'h3 == rs1 ? io_now_reg_3 : _GEN_2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_4 = 5'h4 == rs1 ? io_now_reg_4 : _GEN_3; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5 = 5'h5 == rs1 ? io_now_reg_5 : _GEN_4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_6 = 5'h6 == rs1 ? io_now_reg_6 : _GEN_5; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_7 = 5'h7 == rs1 ? io_now_reg_7 : _GEN_6; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_8 = 5'h8 == rs1 ? io_now_reg_8 : _GEN_7; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_9 = 5'h9 == rs1 ? io_now_reg_9 : _GEN_8; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_10 = 5'ha == rs1 ? io_now_reg_10 : _GEN_9; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_11 = 5'hb == rs1 ? io_now_reg_11 : _GEN_10; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_12 = 5'hc == rs1 ? io_now_reg_12 : _GEN_11; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_13 = 5'hd == rs1 ? io_now_reg_13 : _GEN_12; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_14 = 5'he == rs1 ? io_now_reg_14 : _GEN_13; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_15 = 5'hf == rs1 ? io_now_reg_15 : _GEN_14; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_16 = 5'h10 == rs1 ? io_now_reg_16 : _GEN_15; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_17 = 5'h11 == rs1 ? io_now_reg_17 : _GEN_16; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_18 = 5'h12 == rs1 ? io_now_reg_18 : _GEN_17; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_19 = 5'h13 == rs1 ? io_now_reg_19 : _GEN_18; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_20 = 5'h14 == rs1 ? io_now_reg_20 : _GEN_19; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_21 = 5'h15 == rs1 ? io_now_reg_21 : _GEN_20; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_22 = 5'h16 == rs1 ? io_now_reg_22 : _GEN_21; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_23 = 5'h17 == rs1 ? io_now_reg_23 : _GEN_22; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_24 = 5'h18 == rs1 ? io_now_reg_24 : _GEN_23; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_25 = 5'h19 == rs1 ? io_now_reg_25 : _GEN_24; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_26 = 5'h1a == rs1 ? io_now_reg_26 : _GEN_25; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_27 = 5'h1b == rs1 ? io_now_reg_27 : _GEN_26; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_28 = 5'h1c == rs1 ? io_now_reg_28 : _GEN_27; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_29 = 5'h1d == rs1 ? io_now_reg_29 : _GEN_28; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_30 = 5'h1e == rs1 ? io_now_reg_30 : _GEN_29; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_31 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs1_37 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [11:0] _imm_11_0_T_27 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_26 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_25 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_24 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_23 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_22 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_21 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_20 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_19 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_18 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_17 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_16 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_15 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_14 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_13 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_12 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_11 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_10 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_9 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_8 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_7 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_6 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_5 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_4 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_3 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_2 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_1 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _GEN_65 = _T_1 ? inst[31:20] : 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire [11:0] _GEN_136 = _T_7 ? inst[31:20] : _GEN_65; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_207 = _T_13 ? inst[31:20] : _GEN_136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_278 = _T_19 ? inst[31:20] : _GEN_207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_349 = _T_25 ? inst[31:20] : _GEN_278; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_420 = _T_31 ? inst[31:20] : _GEN_349; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_491 = _T_37 ? inst[31:20] : _GEN_420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_562 = _T_43 ? inst[31:20] : _GEN_491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_633 = _T_49 ? inst[31:20] : _GEN_562; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1735 = _T_157 ? inst[31:20] : _GEN_633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1998 = _T_348 ? inst[31:20] : _GEN_1735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2111 = _T_368 ? inst[31:20] : _GEN_1998; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2224 = _T_388 ? inst[31:20] : _GEN_2111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2302 = _T_408 ? inst[31:20] : _GEN_2224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2415 = _T_427 ? inst[31:20] : _GEN_2302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2515 = _T_518 ? inst[31:20] : _GEN_2415; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2533 = _T_524 ? inst[31:20] : _GEN_2515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2544 = _T_533 ? inst[31:20] : _GEN_2533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4912 = _T_868 ? inst[31:20] : _GEN_2544; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4933 = _T_875 ? inst[31:20] : _GEN_4912; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4947 = _T_882 ? inst[31:20] : _GEN_4933; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4954 = _T_888 ? inst[31:20] : _GEN_4947; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5097 = _T_894 ? inst[31:20] : _GEN_4954; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5269 = _T_927 ? inst[31:20] : _GEN_5097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5441 = _T_967 ? inst[31:20] : _GEN_5269; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5629 = _T_1007 ? inst[31:20] : _GEN_5441; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5801 = _T_1041 ? inst[31:20] : _GEN_5629; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5973 = _T_1082 ? inst[31:20] : _GEN_5801; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] imm_11_0 = io_valid ? _GEN_5973 : 12'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire [11:0] _GEN_6105 = imm_11_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire  imm_signBit_45 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_258 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_259 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_260 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_44 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_255 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_256 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_257 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_43 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_252 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_253 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_254 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_42 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_249 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_250 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_251 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_41 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_246 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_247 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_248 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_40 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_243 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_244 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_245 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_39 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_240 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_241 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_242 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_38 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_237 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_238 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_239 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_37 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_234 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_235 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_236 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_36 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_231 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_232 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_233 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_740 = inst & 32'hec03; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_741 = 32'h8801 == _T_740; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_221 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_222 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_hi_hi_19 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_223 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_hi_19 = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_224 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_225 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_lo_hi_10 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_226 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_lo_19 = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [5:0] _imm_T_227 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  imm_signBit_35 = _imm_T_227[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_228 = imm_signBit_35; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [25:0] _imm_T_229 = imm_signBit_35 ? 26'h3ffffff : 26'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_230 = {_imm_T_229,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_724 = inst & 32'hec03; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_725 = 32'h8401 == _T_740; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_726 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 15:22]
  wire  _T_727 = ~inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 15:27]
  wire  _T_728 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:19]
  wire [4:0] _T_729 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:29]
  wire [5:0] _T_730 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:14]
  wire  _T_731 = _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:37]
  wire  _T_732 = _T_695 & _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:8]
  wire  _T_733 = 32'h8401 == _T_740 & _T_700; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _imm_T_214 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_215 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_hi_hi_18 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_216 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_hi_18 = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_217 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_218 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_lo_hi_9 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_219 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_lo_18 = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [5:0] _imm_T_220 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [31:0] _T_708 = inst & 32'hec03; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_709 = 32'h8001 == _T_740; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_710 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 15:22]
  wire  _T_711 = ~inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 15:27]
  wire  _T_712 = inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:19]
  wire [4:0] _T_713 = inst[6:2]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:29]
  wire [5:0] _T_714 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:14]
  wire  _T_715 = _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:37]
  wire  _T_716 = _T_695 & _T_698 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:8]
  wire  _T_717 = 32'h8001 == _T_740 & _T_700; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _imm_T_207 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_208 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_hi_hi_17 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_209 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_hi_17 = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_210 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_211 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_lo_hi_8 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_212 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_lo_17 = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [5:0] _imm_T_213 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_200 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_201 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_hi_hi_16 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_202 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_hi_16 = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_203 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_204 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_lo_hi_7 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_205 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_lo_16 = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [5:0] _imm_T_206 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_190 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_191 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_hi_hi_15 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_192 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_hi_15 = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_193 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _imm_T_194 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] imm_lo_hi_6 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  _imm_T_195 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [2:0] imm_lo_15 = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [5:0] _imm_T_196 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  imm_signBit_34 = _imm_T_227[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_197 = imm_signBit_35; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [25:0] _imm_T_198 = imm_signBit_35 ? 26'h3ffffff : 26'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_199 = {_imm_T_229,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_616 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_617 = 32'he001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_177 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_178 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_14 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_179 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_180 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_lo_3 = {inst[5],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [3:0] imm_hi_14 = {inst[12],inst[6],inst[5],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_181 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_182 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_hi_5 = {inst[11],inst[10]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_183 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_184 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_lo_3 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [3:0] imm_lo_14 = {inst[11],inst[10],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [7:0] _imm_T_185 = {inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [8:0] _imm_T_186 = {inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_33 = _imm_T_186[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_187 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [22:0] _imm_T_188 = imm_signBit_33 ? 23'h7fffff : 23'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_189 = {_imm_T_188,inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_607 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_608 = 32'hc001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_164 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_165 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_13 = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_166 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_167 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_lo_2 = {inst[5],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [3:0] imm_hi_13 = {inst[12],inst[6],inst[5],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_168 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_169 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_hi_4 = {inst[11],inst[10]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_170 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_171 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_lo_2 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [3:0] imm_lo_13 = {inst[11],inst[10],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [7:0] _imm_T_172 = {inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [8:0] _imm_T_173 = {inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_32 = _imm_T_186[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_174 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [22:0] _imm_T_175 = imm_signBit_33 ? 23'h7fffff : 23'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_176 = {_imm_T_188,inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_583 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_584 = 32'h2001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_585 = 32'h2001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _imm_T_148 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_149 = inst[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_hi_1 = {inst[12],inst[8]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_150 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_hi_12 = {inst[12],inst[8],inst[10]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_151 = inst[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_152 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_lo_hi_1 = {inst[9],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_153 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_lo_1 = {inst[9],inst[6],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [5:0] imm_hi_12 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_154 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_155 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_hi_hi_1 = {inst[2],inst[11]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_156 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_lo_hi_3 = {inst[2],inst[11],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_157 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_158 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_lo_1 = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [4:0] imm_lo_12 = {inst[2],inst[11],inst[5],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [10:0] _imm_T_159 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [11:0] _imm_T_160 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_31 = _imm_T_160[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_161 = imm_signBit_31; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_162 = imm_signBit_31 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_163 = {_imm_T_162,inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_578 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_579 = 32'ha001 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_132 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_133 = inst[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_hi = {inst[12],inst[8]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_134 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_hi_11 = {inst[12],inst[8],inst[10]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_135 = inst[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_136 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_lo_hi = {inst[9],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_137 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_lo = {inst[9],inst[6],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [5:0] imm_hi_11 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_138 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_139 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_hi_hi = {inst[2],inst[11]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_140 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_lo_hi_2 = {inst[2],inst[11],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_141 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_142 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_lo = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [4:0] imm_lo_11 = {inst[2],inst[11],inst[5],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [10:0] _imm_T_143 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [11:0] _imm_T_144 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_30 = _imm_T_160[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_145 = imm_signBit_31; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_146 = imm_signBit_31 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_147 = {_imm_T_162,inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_566 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_567 = 32'hc000 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_124 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_125 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_10 = {inst[5],inst[12]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_126 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_10 = {inst[5],inst[12],inst[11]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_127 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_128 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_10 = {inst[10],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [4:0] _imm_T_129 = {inst[5],inst[12],inst[11],inst[10],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [6:0] _imm_T_130 = {inst[5],inst[12],inst[11],inst[10],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire [31:0] _imm_T_131 = {25'h0,inst[5],inst[12],inst[11],inst[10],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _T_557 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_558 = 32'h4000 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_116 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_117 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_9 = {inst[5],inst[12]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_118 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_9 = {inst[5],inst[12],inst[11]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_119 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_120 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_9 = {inst[10],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [4:0] _imm_T_121 = {inst[5],inst[12],inst[11],inst[10],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [6:0] _imm_T_122 = {inst[5],inst[12],inst[11],inst[10],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire [31:0] _imm_T_123 = {25'h0,inst[5],inst[12],inst[11],inst[10],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _T_548 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_549 = 32'hc002 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _imm_T_107 = inst[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_108 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_8 = {inst[8],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_109 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_8 = {inst[8],inst[7],inst[12]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_110 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_111 = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_hi_1 = {inst[11],inst[10]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_112 = inst[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_lo_8 = {inst[11],inst[10],inst[9]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [5:0] _imm_T_113 = {inst[8],inst[7],inst[12],inst[11],inst[10],inst[9]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [7:0] _imm_T_114 = {inst[8],inst[7],inst[12],inst[11],inst[10],inst[9],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire [31:0] _imm_T_115 = {24'h0,inst[8],inst[7],inst[12],inst[11],inst[10],inst[9],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  _imm_T_98 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_99 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_hi_hi_7 = {inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_100 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_hi_7 = {inst[3],inst[2],inst[12]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_101 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _imm_T_102 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] imm_lo_hi = {inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire  _imm_T_103 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [2:0] imm_lo_7 = {inst[6],inst[5],inst[4]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [5:0] _imm_T_104 = {inst[3],inst[2],inst[12],inst[6],inst[5],inst[4]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [7:0] _imm_T_105 = {inst[3],inst[2],inst[12],inst[6],inst[5],inst[4],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire [31:0] _imm_T_106 = {24'h0,inst[3],inst[2],inst[12],inst[6],inst[5],inst[4],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  imm_signBit_29 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_95 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_96 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_97 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_28 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_92 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_93 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_94 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_27 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_89 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_90 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_91 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [6:0] _imm_11_5_T_2 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _imm_11_5_T_1 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _imm_11_5_T = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _GEN_2461 = _T_447 ? inst[31:25] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [6:0] _GEN_2481 = _T_470 ? inst[31:25] : _GEN_2461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2501 = _T_494 ? inst[31:25] : _GEN_2481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] imm_11_5 = io_valid ? _GEN_2501 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [6:0] _GEN_6162 = imm_11_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [14:0] _T_497 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_498 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _imm_4_0_T_2 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_473 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_474 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _imm_4_0_T_1 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_450 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_451 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _imm_4_0_T = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_2465 = _T_447 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [4:0] _GEN_2485 = _T_470 ? inst[11:7] : _GEN_2465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2505 = _T_494 ? inst[11:7] : _GEN_2485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] imm_4_0 = io_valid ? _GEN_2505 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [4:0] _GEN_6163 = imm_4_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [11:0] _imm_T_85 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_26 = _imm_T_85[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_86 = imm_signBit_26; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_87 = imm_signBit_26 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_88 = {_imm_T_87,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [11:0] _imm_T_81 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_25 = _imm_T_85[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_82 = imm_signBit_26; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_83 = imm_signBit_26 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_84 = {_imm_T_87,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [11:0] _imm_T_77 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_24 = _imm_T_85[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_78 = imm_signBit_26; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_79 = imm_signBit_26 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_80 = {_imm_T_87,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_23 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_74 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_75 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_76 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_22 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_71 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_72 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_73 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_21 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_68 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_69 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_70 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_20 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_65 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_66 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_67 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_19 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_62 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_63 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_64 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _imm_12_T_5 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_4 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_3 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_2 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_1 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _GEN_1789 = _T_182 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire  _GEN_1814 = _T_209 ? inst[31] : _GEN_1789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1839 = _T_236 ? inst[31] : _GEN_1814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1864 = _T_265 ? inst[31] : _GEN_1839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1889 = _T_292 ? inst[31] : _GEN_1864; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1914 = _T_321 ? inst[31] : _GEN_1889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_12 = io_valid & _GEN_1914; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire  _GEN_6155 = imm_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire [14:0] _T_325 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_326 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_327 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_6 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_296 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_297 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_298 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_5 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_269 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_270 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_271 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_4 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_240 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_241 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_242 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_3 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_213 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_214 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_215 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_2 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_186 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_187 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_188 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_1 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_132 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_133 = 32'h6f == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_134 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [20:0] _T_135 = inst[20:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T = inst[20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _GEN_1623 = _T_133 & inst[20]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire  _GEN_1795 = _T_182 ? inst[7] : _GEN_1623; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1820 = _T_209 ? inst[7] : _GEN_1795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1845 = _T_236 ? inst[7] : _GEN_1820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1870 = _T_265 ? inst[7] : _GEN_1845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1895 = _T_292 ? inst[7] : _GEN_1870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1920 = _T_321 ? inst[7] : _GEN_1895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_11 = io_valid & _GEN_1920; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire  _GEN_6148 = imm_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire [1:0] imm_hi_hi_6 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [5:0] _imm_10_5_T_5 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_4 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_3 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_2 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_1 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _GEN_1790 = _T_182 ? inst[30:25] : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [5:0] _GEN_1815 = _T_209 ? inst[30:25] : _GEN_1790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1840 = _T_236 ? inst[30:25] : _GEN_1815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1865 = _T_265 ? inst[30:25] : _GEN_1840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1890 = _T_292 ? inst[30:25] : _GEN_1865; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1915 = _T_321 ? inst[30:25] : _GEN_1890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] imm_10_5 = io_valid ? _GEN_1915 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [5:0] _GEN_6156 = imm_10_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [7:0] imm_hi_6 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [3:0] _imm_4_1_T_5 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_4 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_3 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_2 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_1 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _GEN_1794 = _T_182 ? inst[11:8] : 4'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [3:0] _GEN_1819 = _T_209 ? inst[11:8] : _GEN_1794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1844 = _T_236 ? inst[11:8] : _GEN_1819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1869 = _T_265 ? inst[11:8] : _GEN_1844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1894 = _T_292 ? inst[11:8] : _GEN_1869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1919 = _T_321 ? inst[11:8] : _GEN_1894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] imm_4_1 = io_valid ? _GEN_1919 : 4'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [3:0] _GEN_6157 = imm_4_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [4:0] imm_lo_6 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_58 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_18 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_59 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_60 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_61 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_5 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_5 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_5 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_54 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_17 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_55 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_56 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_57 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_4 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_4 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_4 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_50 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_16 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_51 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_52 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_53 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_3 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_3 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_3 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_46 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_15 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_47 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_48 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_49 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_2 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_2 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_2 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_42 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_14 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_43 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_44 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_45 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_1 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_1 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_1 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_38 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_13 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_39 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_40 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_41 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_12 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_35 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_36 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_37 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _imm_20_T = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _GEN_1621 = _T_133 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire  imm_20 = io_valid & _GEN_1621; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire  _GEN_6146 = imm_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire [19:0] _T_136 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _imm_19_12_T = inst[19:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [7:0] _GEN_1624 = _T_133 ? inst[19:12] : 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [7:0] imm_19_12 = io_valid ? _GEN_1624 : 8'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [7:0] _GEN_6149 = imm_19_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [8:0] imm_hi_hi = {imm_20,imm_19_12}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire [9:0] imm_hi = {imm_20,imm_19_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire [9:0] _imm_10_1_T = inst[30:21]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [9:0] _GEN_1622 = _T_133 ? inst[30:21] : 10'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [9:0] imm_10_1 = io_valid ? _GEN_1622 : 10'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [9:0] _GEN_6147 = imm_10_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [10:0] imm_lo = {imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire [20:0] _imm_T_31 = {imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire  imm_signBit_11 = _imm_T_31[20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_32 = imm_signBit_11; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [10:0] _imm_T_33 = imm_signBit_11 ? 11'h7ff : 11'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_34 = {_imm_T_33,imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_58 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_59 = 32'h17 == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _imm_31_12_T_1 = inst[31:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_54 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_55 = 32'h37 == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _imm_31_12_T = inst[31:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [19:0] _GEN_704 = _T_55 ? inst[31:12] : 20'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [19:0] _GEN_773 = _T_59 ? inst[31:12] : _GEN_704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [19:0] imm_31_12 = io_valid ? _GEN_773 : 20'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [19:0] _GEN_6143 = imm_31_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [31:0] _imm_T_29 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire [31:0] _imm_T_30 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire [31:0] _imm_T_27 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire [31:0] _imm_T_28 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire  imm_signBit_8 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_24 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_25 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_26 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_7 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_21 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_22 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_23 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_6 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_18 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_19 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_20 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_5 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_15 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_16 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_17 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_4 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_12 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_13 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_14 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_3 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_9 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_10 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_11 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_2 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_6 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_7 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_8 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_1 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_3 = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_4 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_5 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T = imm_signBit_45; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_1 = imm_signBit_45 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_2 = {_imm_T_259,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_70 = _T_1 ? _imm_T_260 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 22:24]
  wire [31:0] _GEN_141 = _T_7 ? _imm_T_260 : _GEN_70; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_212 = _T_13 ? _imm_T_260 : _GEN_141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_283 = _T_19 ? _imm_T_260 : _GEN_212; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_354 = _T_25 ? _imm_T_260 : _GEN_283; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_425 = _T_31 ? _imm_T_260 : _GEN_354; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_496 = _T_37 ? _imm_T_260 : _GEN_425; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_567 = _T_43 ? _imm_T_260 : _GEN_496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_638 = _T_49 ? _imm_T_260 : _GEN_567; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_707 = _T_55 ? _imm_T_29 : _GEN_638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [31:0] _GEN_776 = _T_59 ? _imm_T_29 : _GEN_707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [31:0] _GEN_1627 = _T_133 ? _imm_T_34 : _GEN_776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:127]
  wire [31:0] _GEN_1740 = _T_157 ? _imm_T_260 : _GEN_1627; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_1797 = _T_182 ? _imm_T_61 : _GEN_1740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1822 = _T_209 ? _imm_T_61 : _GEN_1797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1847 = _T_236 ? _imm_T_61 : _GEN_1822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1872 = _T_265 ? _imm_T_61 : _GEN_1847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1897 = _T_292 ? _imm_T_61 : _GEN_1872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1922 = _T_321 ? _imm_T_61 : _GEN_1897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_2003 = _T_348 ? _imm_T_260 : _GEN_1922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2116 = _T_368 ? _imm_T_260 : _GEN_2003; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2229 = _T_388 ? _imm_T_260 : _GEN_2116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2307 = _T_408 ? _imm_T_260 : _GEN_2229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2420 = _T_427 ? _imm_T_260 : _GEN_2307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2467 = _T_447 ? _imm_T_88 : _GEN_2420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [31:0] _GEN_2487 = _T_470 ? _imm_T_88 : _GEN_2467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [31:0] _GEN_2507 = _T_494 ? _imm_T_88 : _GEN_2487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [31:0] _GEN_2520 = _T_518 ? _imm_T_260 : _GEN_2507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2538 = _T_524 ? _imm_T_260 : _GEN_2520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2549 = _T_533 ? _imm_T_260 : _GEN_2538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2589 = _T_542 ? _imm_T_106 : _GEN_2549; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 140:20]
  wire [31:0] _GEN_2630 = _T_549 ? _imm_T_115 : _GEN_2589; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 145:11]
  wire [31:0] _GEN_2706 = _T_558 ? _imm_T_131 : _GEN_2630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 151:28]
  wire [31:0] _GEN_2813 = _T_567 ? _imm_T_131 : _GEN_2706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 156:11]
  wire [31:0] _GEN_2822 = _T_579 ? _imm_T_163 : _GEN_2813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 162:25]
  wire [31:0] _GEN_2829 = _T_584 ? _imm_T_163 : _GEN_2822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 168:25]
  wire [31:0] _GEN_2891 = _T_608 ? _imm_T_189 : _GEN_2829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 188:11]
  wire [31:0] _GEN_2935 = _T_617 ? _imm_T_189 : _GEN_2891; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 196:11]
  wire [31:0] _GEN_2977 = _T_629 ? _imm_T_230 : _GEN_2935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 206:20]
  wire [31:0] _GEN_3300 = _T_702 ? {{26'd0}, _imm_T_227} : _GEN_2977; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 232:20]
  wire [31:0] _GEN_3404 = _T_717 ? {{26'd0}, _imm_T_227} : _GEN_3300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 237:28]
  wire [31:0] _GEN_3508 = _T_733 ? {{26'd0}, _imm_T_227} : _GEN_3404; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 242:28]
  wire [31:0] _GEN_3612 = _T_741 ? _imm_T_230 : _GEN_3508; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 247:28]
  wire [31:0] _GEN_4917 = _T_868 ? _imm_T_260 : _GEN_3612; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_4938 = _T_875 ? _imm_T_260 : _GEN_4917; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _GEN_4952 = _T_882 ? _imm_T_260 : _GEN_4938; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28]
  wire [31:0] _GEN_4959 = _T_888 ? _imm_T_260 : _GEN_4952; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28]
  wire [31:0] _GEN_5102 = _T_894 ? _imm_T_260 : _GEN_4959; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5274 = _T_927 ? _imm_T_260 : _GEN_5102; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5446 = _T_967 ? _imm_T_260 : _GEN_5274; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_5634 = _T_1007 ? _imm_T_260 : _GEN_5446; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_5806 = _T_1041 ? _imm_T_260 : _GEN_5634; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_5978 = _T_1082 ? _imm_T_260 : _GEN_5806; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] imm = io_valid ? _GEN_5978 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [31:0] _GEN_6110 = imm; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [32:0] _T_432 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:47]
  wire [31:0] _T_433 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:47]
  wire [2:0] _T_438 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_439 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_442 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_436 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_437 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_440 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_434 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_435 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_441 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_443 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_445 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_423 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [4:0] _rs2_T_31 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_30 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_29 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_28 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_27 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_26 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_25 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_24 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_770 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs2_T_23 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_758 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs2_T_22 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_605 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs2_T_21 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_596 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs2_T_20 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_550 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 114:97]
  wire [12:0] _T_551 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [6:0] _T_552 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs2_T_19 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_18 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_17 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_16 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_15 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_14 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_13 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_12 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_11 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_10 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_9 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_8 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_7 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_6 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_5 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_4 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_3 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_2 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_1 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_875 = _T_63 ? inst[24:20] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [4:0] _GEN_946 = _T_70 ? inst[24:20] : _GEN_875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1017 = _T_77 ? inst[24:20] : _GEN_946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1088 = _T_84 ? inst[24:20] : _GEN_1017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1159 = _T_91 ? inst[24:20] : _GEN_1088; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1230 = _T_98 ? inst[24:20] : _GEN_1159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1301 = _T_105 ? inst[24:20] : _GEN_1230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1372 = _T_112 ? inst[24:20] : _GEN_1301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1443 = _T_119 ? inst[24:20] : _GEN_1372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1514 = _T_126 ? inst[24:20] : _GEN_1443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1791 = _T_182 ? inst[24:20] : _GEN_1514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1816 = _T_209 ? inst[24:20] : _GEN_1791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1841 = _T_236 ? inst[24:20] : _GEN_1816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1866 = _T_265 ? inst[24:20] : _GEN_1841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1891 = _T_292 ? inst[24:20] : _GEN_1866; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1916 = _T_321 ? inst[24:20] : _GEN_1891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2462 = _T_447 ? inst[24:20] : _GEN_1916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2482 = _T_470 ? inst[24:20] : _GEN_2462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2502 = _T_494 ? inst[24:20] : _GEN_2482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2628 = _T_549 ? inst[6:2] : _GEN_2502; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2836 = _T_593 ? inst[6:2] : _GEN_2628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2844 = _T_602 ? inst[6:2] : _GEN_2836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3680 = _T_755 ? inst[6:2] : _GEN_2844; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3750 = _T_767 ? inst[6:2] : _GEN_3680; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4366 = _T_812 ? inst[24:20] : _GEN_3750; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4437 = _T_819 ? inst[24:20] : _GEN_4366; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4508 = _T_826 ? inst[24:20] : _GEN_4437; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4579 = _T_833 ? inst[24:20] : _GEN_4508; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4650 = _T_840 ? inst[24:20] : _GEN_4579; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4721 = _T_847 ? inst[24:20] : _GEN_4650; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4792 = _T_854 ? inst[24:20] : _GEN_4721; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4863 = _T_861 ? inst[24:20] : _GEN_4792; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs2 = io_valid ? _GEN_4863 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [4:0] _GEN_6145 = rs2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [2:0] _T_417 = rs2[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_418 = rs2[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_421 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_415 = rs2[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_416 = rs2[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_419 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_413 = rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_414 = ~rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_420 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_422 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_424 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_425 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 107:10]
  wire  _T_405 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_33 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_393 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:47]
  wire [31:0] _T_394 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:47]
  wire [2:0] _T_399 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_400 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_403 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_397 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_398 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_401 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_395 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_396 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_402 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_404 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_406 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_385 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_30 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_373 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:47]
  wire [31:0] _T_374 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:47]
  wire [2:0] _T_379 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_380 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_383 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_377 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_378 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_381 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_375 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_376 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_382 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_384 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_386 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_365 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_27 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_353 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:47]
  wire [31:0] _T_354 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:47]
  wire [2:0] _T_359 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_360 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_363 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_357 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_358 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_361 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_355 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_356 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_362 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_364 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_366 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _exceptionVec_WIRE_4 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_1995 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_2039 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2108 = _T_435 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2152 = _T_368 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2221 = _T_437 ? _GEN_2152 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2265 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2267 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2308 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2412 = _T_435 ? _GEN_2265 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2456 = _T_427 ? _GEN_2412 : _GEN_2265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  exceptionVec_4 = io_valid & _GEN_2456; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6161 = exceptionVec_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_4 = exceptionVec_4 ? 5'h4 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _T_512 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_44 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_500 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:47]
  wire [31:0] _T_501 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:47]
  wire [2:0] _T_506 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_507 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_510 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_504 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_505 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_508 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_502 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_503 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_509 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_511 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_513 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_488 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_41 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_476 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:47]
  wire [31:0] _T_477 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:47]
  wire [2:0] _T_482 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_483 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_486 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_480 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_481 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_484 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_478 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_479 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_485 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_487 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_489 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_463 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [2:0] _T_457 = rs2[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_458 = rs2[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_461 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_455 = rs2[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_456 = rs2[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_459 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_453 = rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_454 = ~rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_460 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_462 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_464 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_465 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 107:10]
  wire  _exceptionVec_WIRE_6 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2458 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 107:36 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_2468 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2478 = _T_435 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2492 = _T_470 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2498 = _T_437 ? _GEN_2492 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2512 = _T_494 ? _GEN_2498 : _GEN_2492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  exceptionVec_6 = io_valid & _GEN_2512; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6164 = exceptionVec_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_5 = exceptionVec_6 ? 5'h6 : _exceptionNO_T_4; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [1:0] now_internal_privilegeMode = io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_529 = 2'h3 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _exceptionVec_WIRE_8 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _T_530 = 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _T_531 = 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2523 = 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2527 = 2'h1 == io_now_internal_privilegeMode ? 1'h0 : 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2531 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : _GEN_2527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2542 = _T_524 & _GEN_2531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_8 = io_valid & _GEN_2542; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6172 = exceptionVec_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_6 = exceptionVec_8 ? 5'h8 : _exceptionNO_T_5; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_9 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2525 = 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2530 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2541 = _T_524 & _GEN_2530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_9 = io_valid & _GEN_2541; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6171 = exceptionVec_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_7 = exceptionVec_9 ? 5'h9 : _exceptionNO_T_6; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_11 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2528 = 2'h3 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2539 = _T_524 & _T_529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_11 = io_valid & _GEN_2539; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6170 = exceptionVec_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_8 = exceptionVec_11 ? 5'hb : _exceptionNO_T_7; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _now_reg_rs1_26 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_809 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_810 = 5'h1 == rs2 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_811 = 5'h2 == rs2 ? io_now_reg_2 : _GEN_810; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_812 = 5'h3 == rs2 ? io_now_reg_3 : _GEN_811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_813 = 5'h4 == rs2 ? io_now_reg_4 : _GEN_812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_814 = 5'h5 == rs2 ? io_now_reg_5 : _GEN_813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_815 = 5'h6 == rs2 ? io_now_reg_6 : _GEN_814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_816 = 5'h7 == rs2 ? io_now_reg_7 : _GEN_815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_817 = 5'h8 == rs2 ? io_now_reg_8 : _GEN_816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_818 = 5'h9 == rs2 ? io_now_reg_9 : _GEN_817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_819 = 5'ha == rs2 ? io_now_reg_10 : _GEN_818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_820 = 5'hb == rs2 ? io_now_reg_11 : _GEN_819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_821 = 5'hc == rs2 ? io_now_reg_12 : _GEN_820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_822 = 5'hd == rs2 ? io_now_reg_13 : _GEN_821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_823 = 5'he == rs2 ? io_now_reg_14 : _GEN_822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_824 = 5'hf == rs2 ? io_now_reg_15 : _GEN_823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_825 = 5'h10 == rs2 ? io_now_reg_16 : _GEN_824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_826 = 5'h11 == rs2 ? io_now_reg_17 : _GEN_825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_827 = 5'h12 == rs2 ? io_now_reg_18 : _GEN_826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_828 = 5'h13 == rs2 ? io_now_reg_19 : _GEN_827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_829 = 5'h14 == rs2 ? io_now_reg_20 : _GEN_828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_830 = 5'h15 == rs2 ? io_now_reg_21 : _GEN_829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_831 = 5'h16 == rs2 ? io_now_reg_22 : _GEN_830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_832 = 5'h17 == rs2 ? io_now_reg_23 : _GEN_831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_833 = 5'h18 == rs2 ? io_now_reg_24 : _GEN_832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_834 = 5'h19 == rs2 ? io_now_reg_25 : _GEN_833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_835 = 5'h1a == rs2 ? io_now_reg_26 : _GEN_834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_836 = 5'h1b == rs2 ? io_now_reg_27 : _GEN_835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_837 = 5'h1c == rs2 ? io_now_reg_28 : _GEN_836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_838 = 5'h1d == rs2 ? io_now_reg_29 : _GEN_837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_839 = 5'h1e == rs2 ? io_now_reg_30 : _GEN_838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_840 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _now_reg_rs2_14 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_329 = _GEN_31 >= _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:25]
  wire [31:0] now_csr_misa = io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_330 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_331 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_332 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_345 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] now_pc = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [32:0] _T_333 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:49]
  wire [31:0] _T_334 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:49]
  wire [2:0] _T_339 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_340 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_343 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_337 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_338 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_341 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_335 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_336 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_342 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_344 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_346 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_25 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _T_300 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:25]
  wire [31:0] _now_reg_rs2_13 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_301 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:48]
  wire  _T_302 = $signed(_T_300) >= $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:32]
  wire  _T_303 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_304 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_305 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_318 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_306 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:49]
  wire [31:0] _T_307 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:49]
  wire [2:0] _T_312 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_313 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_316 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_310 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_311 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_314 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_308 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_309 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_315 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_317 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_319 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_24 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_12 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_273 = _GEN_31 < _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:25]
  wire  _T_274 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_275 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_276 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_289 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_277 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:49]
  wire [31:0] _T_278 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:49]
  wire [2:0] _T_283 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_284 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_287 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_281 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_282 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_285 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_279 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_280 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_286 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_288 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_290 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_23 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _T_244 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:25]
  wire [31:0] _now_reg_rs2_11 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_245 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:47]
  wire  _T_246 = $signed(_T_300) < $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:32]
  wire  _T_247 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_248 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_249 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_262 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_250 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:49]
  wire [31:0] _T_251 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:49]
  wire [2:0] _T_256 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_257 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_260 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_254 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_255 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_258 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_252 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_253 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_259 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_261 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_263 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_22 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_10 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_217 = _GEN_31 != _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:25]
  wire  _T_218 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_219 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_220 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_233 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_221 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:49]
  wire [31:0] _T_222 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:49]
  wire [2:0] _T_227 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_228 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_231 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_225 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_226 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_229 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_223 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_224 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_230 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_232 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_234 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_21 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_9 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_190 = _GEN_31 == _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:25]
  wire  _T_191 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_192 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_193 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_206 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_194 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:49]
  wire [31:0] _T_195 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:49]
  wire [2:0] _T_200 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_201 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_204 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_198 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_199 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_202 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_196 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_197 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_203 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_205 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_207 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_162 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_163 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_164 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_179 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_18 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_165 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:58]
  wire [31:0] _T_166 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:58]
  wire [30:0] _T_167 = _T_433[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:64]
  wire [31:0] _T_168 = {_T_433[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:43]
  wire [2:0] _T_173 = _T_168[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_174 = _T_168[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_177 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_171 = _T_168[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_172 = _T_168[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_175 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_169 = _T_168[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_170 = ~_T_168[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_176 = 2'h1 == _T_332 ? _T_170 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_178 = 2'h2 == _T_332 ? _T_172 : _T_176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_180 = 2'h3 == _T_332 ? _T_174 : _T_178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_139 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_140 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_141 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_154 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_142 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:47]
  wire [31:0] _T_143 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:47]
  wire [2:0] _T_148 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_149 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_152 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_146 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_147 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_150 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_144 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_145 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_151 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_153 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_155 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _exceptionVec_WIRE_0 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_1618 = _T_346 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_1663 = _T_133 & _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_1732 = _T_180 ? _GEN_1663 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1776 = _T_157 ? _GEN_1732 : _GEN_1663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1781 = _T_346 ? _GEN_1776 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1786 = _GEN_31 == _GEN_840 ? _GEN_1781 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1801 = _T_182 ? _GEN_1786 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1806 = _T_346 ? _GEN_1801 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1811 = _GEN_31 != _GEN_840 ? _GEN_1806 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1826 = _T_209 ? _GEN_1811 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1831 = _T_346 ? _GEN_1826 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1836 = $signed(_T_300) < $signed(_T_301) ? _GEN_1831 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1851 = _T_236 ? _GEN_1836 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1856 = _T_346 ? _GEN_1851 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1861 = _GEN_31 < _GEN_840 ? _GEN_1856 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1876 = _T_265 ? _GEN_1861 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1881 = _T_346 ? _GEN_1876 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1886 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1881 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1901 = _T_292 ? _GEN_1886 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1906 = _T_346 ? _GEN_1901 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1911 = _GEN_31 >= _GEN_840 ? _GEN_1906 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1926 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  exceptionVec_0 = io_valid & _GEN_1926; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6153 = exceptionVec_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_9 = exceptionVec_0 ? 5'h0 : _exceptionNO_T_8; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _T_796 = inst & 32'hfc63; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_797 = 32'h8c01 == _T_796; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_788 = inst & 32'hfc63; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_789 = 32'h8c21 == _T_796; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_780 = inst & 32'hfc63; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_781 = 32'h8c41 == _T_796; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_772 = inst & 32'hfc63; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_773 = 32'h8c61 == _T_796; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_680 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_681 = 32'h0 == _T_690; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire [7:0] _T_682 = inst[12:5]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 23:88]
  wire  _T_683 = inst[12:5] != 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 23:96]
  wire  _T_684 = 32'h0 == _T_690 & _T_683; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _GEN_64 = _T_1 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 125:24 128:24]
  wire  _GEN_135 = _T_7 ? 1'h0 : _GEN_64; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_206 = _T_13 ? 1'h0 : _GEN_135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_277 = _T_19 ? 1'h0 : _GEN_206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_348 = _T_25 ? 1'h0 : _GEN_277; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_419 = _T_31 ? 1'h0 : _GEN_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_490 = _T_37 ? 1'h0 : _GEN_419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_561 = _T_43 ? 1'h0 : _GEN_490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_632 = _T_49 ? 1'h0 : _GEN_561; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_703 = _T_55 ? 1'h0 : _GEN_632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_772 = _T_59 ? 1'h0 : _GEN_703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_873 = _T_63 ? 1'h0 : _GEN_772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_944 = _T_70 ? 1'h0 : _GEN_873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1015 = _T_77 ? 1'h0 : _GEN_944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1086 = _T_84 ? 1'h0 : _GEN_1015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1157 = _T_91 ? 1'h0 : _GEN_1086; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1228 = _T_98 ? 1'h0 : _GEN_1157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1299 = _T_105 ? 1'h0 : _GEN_1228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1370 = _T_112 ? 1'h0 : _GEN_1299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1441 = _T_119 ? 1'h0 : _GEN_1370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1512 = _T_126 ? 1'h0 : _GEN_1441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1620 = _T_133 ? 1'h0 : _GEN_1512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1734 = _T_157 ? 1'h0 : _GEN_1620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1788 = _T_182 ? 1'h0 : _GEN_1734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1813 = _T_209 ? 1'h0 : _GEN_1788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1838 = _T_236 ? 1'h0 : _GEN_1813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1863 = _T_265 ? 1'h0 : _GEN_1838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1888 = _T_292 ? 1'h0 : _GEN_1863; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1913 = _T_321 ? 1'h0 : _GEN_1888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1997 = _T_348 ? 1'h0 : _GEN_1913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2110 = _T_368 ? 1'h0 : _GEN_1997; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2223 = _T_388 ? 1'h0 : _GEN_2110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2301 = _T_408 ? 1'h0 : _GEN_2223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2414 = _T_427 ? 1'h0 : _GEN_2301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2460 = _T_447 ? 1'h0 : _GEN_2414; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2480 = _T_470 ? 1'h0 : _GEN_2460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2500 = _T_494 ? 1'h0 : _GEN_2480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2514 = _T_518 ? 1'h0 : _GEN_2500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2532 = _T_524 ? 1'h0 : _GEN_2514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2543 = _T_533 ? 1'h0 : _GEN_2532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2582 = _T_542 ? 1'h0 : _GEN_2543; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2625 = _T_549 ? 1'h0 : _GEN_2582; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2699 = _T_558 ? 1'h0 : _GEN_2625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2806 = _T_567 ? 1'h0 : _GEN_2699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2818 = _T_579 ? 1'h0 : _GEN_2806; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2825 = _T_584 ? 1'h0 : _GEN_2818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2833 = _T_593 ? 1'h0 : _GEN_2825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2841 = _T_602 ? 1'h0 : _GEN_2833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2884 = _T_608 ? 1'h0 : _GEN_2841; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2928 = _T_617 ? 1'h0 : _GEN_2884; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2970 = _T_629 ? 1'h0 : _GEN_2928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3042 = _T_647 ? 1'h0 : _GEN_2970; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3145 = _T_662 ? 1'h0 : _GEN_3042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3184 = _T_674 ? 1'h0 : _GEN_3145; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3224 = _T_684 ? 1'h0 : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3293 = _T_702 ? 1'h0 : _GEN_3224; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3397 = _T_717 ? 1'h0 : _GEN_3293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3501 = _T_733 ? 1'h0 : _GEN_3397; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3605 = _T_741 ? 1'h0 : _GEN_3501; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3677 = _T_755 ? 1'h0 : _GEN_3605; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3747 = _T_767 ? 1'h0 : _GEN_3677; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3881 = _T_773 ? 1'h0 : _GEN_3747; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4016 = _T_781 ? 1'h0 : _GEN_3881; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4151 = _T_789 ? 1'h0 : _GEN_4016; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4286 = _T_797 ? 1'h0 : _GEN_4151; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4325 = _T_805 ? 1'h0 : _GEN_4286; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4364 = _T_812 ? 1'h0 : _GEN_4325; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4435 = _T_819 ? 1'h0 : _GEN_4364; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4506 = _T_826 ? 1'h0 : _GEN_4435; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4577 = _T_833 ? 1'h0 : _GEN_4506; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4648 = _T_840 ? 1'h0 : _GEN_4577; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4719 = _T_847 ? 1'h0 : _GEN_4648; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4790 = _T_854 ? 1'h0 : _GEN_4719; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4861 = _T_861 ? 1'h0 : _GEN_4790; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4911 = _T_868 ? 1'h0 : _GEN_4861; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4932 = _T_875 ? 1'h0 : _GEN_4911; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4946 = _T_882 ? 1'h0 : _GEN_4932; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4953 = _T_888 ? 1'h0 : _GEN_4946; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5096 = _T_894 ? 1'h0 : _GEN_4953; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5268 = _T_927 ? 1'h0 : _GEN_5096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5440 = _T_967 ? 1'h0 : _GEN_5268; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5628 = _T_1007 ? 1'h0 : _GEN_5440; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5800 = _T_1041 ? 1'h0 : _GEN_5628; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5972 = _T_1082 ? 1'h0 : _GEN_5800; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  illegalInstruction = io_valid & _GEN_5972; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 119:36]
  wire  _GEN_6102 = illegalInstruction; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 119:36]
  wire [11:0] _csrAddr_T_5 = imm[11:0]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:19]
  wire [11:0] _csrAddr_T_4 = imm[11:0]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:19]
  wire [11:0] _csrAddr_T_3 = imm[11:0]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:19]
  wire [11:0] _csrAddr_T_2 = imm[11:0]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:19]
  wire [11:0] _csrAddr_T_1 = imm[11:0]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:19]
  wire [11:0] _csrAddr_T = imm[11:0]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:19]
  wire [11:0] _GEN_5103 = _T_894 ? imm[11:0] : 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:13 82:23 53:25]
  wire [11:0] _GEN_5275 = _T_927 ? imm[11:0] : _GEN_5103; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:13 93:23]
  wire [11:0] _GEN_5447 = _T_967 ? imm[11:0] : _GEN_5275; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 56:13]
  wire [11:0] _GEN_5635 = _T_1007 ? imm[11:0] : _GEN_5447; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 56:13]
  wire [11:0] _GEN_5807 = _T_1041 ? imm[11:0] : _GEN_5635; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 56:13]
  wire [11:0] _GEN_5979 = _T_1082 ? imm[11:0] : _GEN_5807; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 56:13]
  wire [11:0] csrAddr = io_valid ? _GEN_5979 : 12'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 53:25]
  wire [11:0] _GEN_6191 = csrAddr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 53:25]
  wire [1:0] _isIllegalWrite_T_15 = csrAddr[11:10]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:30]
  wire  isIllegalWrite_5 = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _isIllegalWrite_T_17 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:55]
  wire  _isIllegalWrite_T_16 = isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _T_1089 = ~isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:12]
  wire  _T_1090 = rs1 != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:18]
  wire  _has_T_431 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_429 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_427 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_425 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_423 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_421 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_419 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_417 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_415 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_413 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_411 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_409 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_407 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_405 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_406 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_408 = 12'hf11 == csrAddr | 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_410 = 12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_412 = 12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_414 = 12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 ==
    csrAddr))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_416 = 12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr)))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_418 = 12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_420 = 12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_422 = 12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_424 = 12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 ==
    csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr
    )))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_426 = 12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 ==
    csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_428 = 12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 ==
    csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_430 = 12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 ==
    csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_15 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire [1:0] _isIllegalMode_T_5 = csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:59]
  wire  isIllegalMode_5 = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess_5 = isIllegalMode_5 | isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _has_T_377 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_375 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_373 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_371 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_369 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_367 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_365 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_363 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_361 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_359 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_357 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_355 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_353 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_351 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_352 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_354 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_356 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_358 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_360 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_362 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_364 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_366 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_368 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_370 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_372 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_374 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_376 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  has_13 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _T_1087 = ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:29]
  wire  _T_1088 = isIllegalAccess_5 | ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:26]
  wire [1:0] _isIllegalWrite_T_12 = csrAddr[11:10]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:30]
  wire  _isIllegalWrite_T_13 = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire [31:0] _now_reg_rs1_74 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _T_1046 = _GEN_31 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:39]
  wire  _isIllegalWrite_T_14 = ~_T_1046; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:55]
  wire  isIllegalWrite_4 = isIllegalWrite_5 & ~_T_1046; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:51]
  wire  _T_1049 = ~isIllegalWrite_4; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:12]
  wire  _T_1050 = rs1 != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:18]
  wire  _has_T_350 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_348 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_346 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_344 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_342 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_340 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_338 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_336 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_334 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_332 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_330 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_328 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_326 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_324 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_325 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_327 = 12'hf11 == csrAddr | 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_329 = 12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_331 = 12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_333 = 12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 ==
    csrAddr))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_335 = 12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr)))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_337 = 12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_339 = 12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_341 = 12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_343 = 12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 ==
    csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr
    )))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_345 = 12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 ==
    csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_347 = 12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 ==
    csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_349 = 12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 ==
    csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_12 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire [1:0] _isIllegalMode_T_4 = csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:59]
  wire  isIllegalMode_4 = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess_4 = isIllegalMode_5 | isIllegalWrite_4; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _has_T_296 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_294 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_292 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_290 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_288 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_286 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_284 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_282 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_280 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_278 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_276 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_274 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_272 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_270 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_271 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_273 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_275 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_277 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_279 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_281 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_283 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_285 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_287 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_289 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_291 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_293 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_295 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  has_10 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _T_1047 = ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:29]
  wire  _T_1048 = isIllegalAccess_4 | ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:26]
  wire [1:0] _isIllegalWrite_T_9 = csrAddr[11:10]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:30]
  wire  isIllegalWrite_3 = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _isIllegalWrite_T_11 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:55]
  wire  _isIllegalWrite_T_10 = isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _T_1014 = ~isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:12]
  wire  _has_T_269 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_267 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_265 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_263 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_261 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_259 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_257 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_255 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_253 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_251 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_249 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_247 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_245 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_243 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_244 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_246 = 12'hf11 == csrAddr | 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_248 = 12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_250 = 12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_252 = 12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 ==
    csrAddr))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_254 = 12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr)))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_256 = 12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_258 = 12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_260 = 12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_262 = 12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 ==
    csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr
    )))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_264 = 12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 ==
    csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_266 = 12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 ==
    csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_268 = 12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 ==
    csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_9 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire [1:0] _isIllegalMode_T_3 = csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:59]
  wire  isIllegalMode_3 = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess_3 = isIllegalMode_5 | isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _has_T_242 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_240 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_238 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_236 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_234 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_232 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_230 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_228 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_226 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_224 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_222 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_220 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_218 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_216 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_217 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_219 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_221 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_223 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_225 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_227 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_229 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_231 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_233 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_235 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_237 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_239 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_241 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  has_8 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _T_1012 = ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:29]
  wire  _T_1013 = isIllegalAccess_5 | ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:26]
  wire [1:0] _isIllegalWrite_T_6 = csrAddr[11:10]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:30]
  wire  isIllegalWrite_2 = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _isIllegalWrite_T_8 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:55]
  wire  _isIllegalWrite_T_7 = isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _T_974 = ~isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:12]
  wire  _T_975 = rs1 != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:18]
  wire  _has_T_215 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_213 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_211 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_209 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_207 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_205 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_203 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_201 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_199 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_197 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_195 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_193 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_191 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_189 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_190 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_192 = 12'hf11 == csrAddr | 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_194 = 12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_196 = 12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_198 = 12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 ==
    csrAddr))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_200 = 12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr)))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_202 = 12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_204 = 12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_206 = 12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_208 = 12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 ==
    csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr
    )))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_210 = 12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 ==
    csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_212 = 12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 ==
    csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_214 = 12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 ==
    csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_7 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire [1:0] _isIllegalMode_T_2 = csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:59]
  wire  isIllegalMode_2 = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess_2 = isIllegalMode_5 | isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _has_T_161 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_159 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_157 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_155 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_153 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_151 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_149 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_147 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_145 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_143 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_141 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_139 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_137 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_135 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_136 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_138 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_140 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_142 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_144 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_146 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_148 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_150 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_152 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_154 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_156 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_158 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_160 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  has_5 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _T_972 = ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:29]
  wire  _T_973 = isIllegalAccess_5 | ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:26]
  wire [1:0] _isIllegalWrite_T_3 = csrAddr[11:10]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:30]
  wire  _isIllegalWrite_T_4 = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire [31:0] _now_reg_rs1_71 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _T_932 = _GEN_31 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:39]
  wire  _isIllegalWrite_T_5 = ~_T_1046; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:55]
  wire  isIllegalWrite_1 = isIllegalWrite_5 & ~_T_1046; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:51]
  wire  _T_935 = ~isIllegalWrite_4; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:12]
  wire  _T_936 = rs1 != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:18]
  wire  _has_T_134 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_132 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_130 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_128 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_126 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_124 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_122 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_120 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_118 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_116 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_114 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_112 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_110 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_108 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_109 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_111 = 12'hf11 == csrAddr | 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_113 = 12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_115 = 12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_117 = 12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 ==
    csrAddr))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_119 = 12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr)))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_121 = 12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_123 = 12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_125 = 12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_127 = 12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 ==
    csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr
    )))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_129 = 12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 ==
    csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_131 = 12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 ==
    csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_133 = 12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 ==
    csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_4 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire [1:0] _isIllegalMode_T_1 = csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:59]
  wire  isIllegalMode_1 = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess_1 = isIllegalMode_5 | isIllegalWrite_4; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _has_T_80 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_78 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_76 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_74 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_72 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_70 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_68 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_66 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_64 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_62 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_60 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_58 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_56 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_54 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_55 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_57 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_59 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_61 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_63 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_65 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_67 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_69 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_71 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_73 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_75 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_77 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_79 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  has_2 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _T_933 = ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:29]
  wire  _T_934 = isIllegalAccess_4 | ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:26]
  wire [1:0] _isIllegalWrite_T = csrAddr[11:10]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:30]
  wire  isIllegalWrite = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _isIllegalWrite_T_2 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:55]
  wire  _isIllegalWrite_T_1 = isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _T_901 = ~isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:12]
  wire  _has_T_53 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_51 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_49 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_47 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_45 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_43 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_41 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_39 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_37 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_35 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_33 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_31 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_29 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_27 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_28 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_30 = 12'hf11 == csrAddr | 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_32 = 12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_34 = 12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_36 = 12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 ==
    csrAddr))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_38 = 12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr)))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_40 = 12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_42 = 12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_44 = 12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_46 = 12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 ==
    csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr
    )))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_48 = 12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 ==
    csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 ==
    csrAddr | 12'h301 == csrAddr))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_50 = 12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 == csrAddr | (12'h305 ==
    csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 == csrAddr | (12'hf12 ==
    csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_52 = 12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 == csrAddr | (12'h306 ==
    csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 == csrAddr | (12'hf13 ==
    csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_1 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire [1:0] _isIllegalMode_T = csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:59]
  wire  isIllegalMode = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess = isIllegalMode_5 | isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _has_T_26 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_24 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_22 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_20 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_18 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_16 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_14 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_12 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_10 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_8 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_6 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_4 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_2 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_1 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_3 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_5 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_7 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_9 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_11 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_13 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_15 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_17 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_19 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_21 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_23 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _has_T_25 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  has = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 75:51]
  wire  _T_899 = ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:29]
  wire  _T_900 = isIllegalAccess_5 | ~has_15; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:26]
  wire  _T_880 = io_now_internal_privilegeMode == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:37]
  wire  illegalSret = io_now_internal_privilegeMode < 2'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 118:55]
  wire  _illegalSModeSret_T = io_now_internal_privilegeMode == 2'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 119:55]
  wire [31:0] now_csr_mstatus = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _mstatusOld_WIRE_1 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusOld_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_18 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _illegalSModeSret_T_1 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  illegalSModeSret = io_now_internal_privilegeMode == 2'h1 & mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 119:65]
  wire  _T_873 = illegalSret | illegalSModeSret; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:22]
  wire  _exceptionVec_WIRE_2 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_4900 = illegalSret | illegalSModeSret; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:22]
  wire  _GEN_4918 = _T_868 & _T_873; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_4930 = io_now_internal_privilegeMode == 2'h3 ? _GEN_4918 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_4944 = _T_875 ? _GEN_4930 : _GEN_4918; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_4960 = isIllegalAccess_5 | ~has_15 | _GEN_4944; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5050 = has_15 ? _GEN_4960 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5094 = _T_1089 ? _GEN_5050 : _GEN_4960; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire  _GEN_5104 = _T_894 ? _GEN_5094 : _GEN_4944; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire  _GEN_5148 = isIllegalAccess_4 | ~has_15 | _GEN_5104; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5210 = has_15 ? _GEN_5148 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5222 = _T_1090 ? _GEN_5210 : _GEN_5148; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire  _GEN_5266 = _T_1049 ? _GEN_5222 : _GEN_5148; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire  _GEN_5276 = _T_927 ? _GEN_5266 : _GEN_5104; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire  _GEN_5320 = isIllegalAccess_5 | ~has_15 | _GEN_5276; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5382 = has_15 ? _GEN_5320 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5394 = _T_1090 ? _GEN_5382 : _GEN_5320; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire  _GEN_5438 = _T_1089 ? _GEN_5394 : _GEN_5320; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire  _GEN_5448 = _T_967 ? _GEN_5438 : _GEN_5276; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire  _GEN_5492 = isIllegalAccess_5 | ~has_15 | _GEN_5448; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5582 = has_15 ? _GEN_5492 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5626 = _T_1089 ? _GEN_5582 : _GEN_5492; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire  _GEN_5636 = _T_1007 ? _GEN_5626 : _GEN_5448; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire  _GEN_5680 = isIllegalAccess_4 | ~has_15 | _GEN_5636; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5742 = has_15 ? _GEN_5680 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5754 = _T_1090 ? _GEN_5742 : _GEN_5680; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire  _GEN_5798 = ~isIllegalWrite_4 ? _GEN_5754 : _GEN_5680; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire  _GEN_5808 = _T_1041 ? _GEN_5798 : _GEN_5636; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire  _GEN_5852 = isIllegalAccess_5 | ~has_15 | _GEN_5808; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5914 = has_15 ? _GEN_5852 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5926 = rs1 != 5'h0 ? _GEN_5914 : _GEN_5852; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire  _GEN_5970 = ~isIllegalWrite_5 ? _GEN_5926 : _GEN_5852; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire  _GEN_5980 = _T_1082 ? _GEN_5970 : _GEN_5808; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire  _GEN_6025 = illegalInstruction | _GEN_5980; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 144:33]
  wire  exceptionVec_2 = io_valid & _GEN_6025; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6187 = exceptionVec_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_10 = exceptionVec_2 ? 5'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_11 = exceptionVec_2 ? 5'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_12 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_12 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_12 = exceptionVec_2 ? 5'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_3 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2521 = 32'h100073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  exceptionVec_3 = io_valid & _T_518; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_6169 = exceptionVec_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] exceptionNO = exceptionVec_3 ? 5'h3 : _exceptionNO_T_10; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] now_csr_cycle = io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [32:0] _next_csr_cycle_T = io_now_csr_cycle + 32'h1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 126:37]
  wire [31:0] _next_csr_cycle_T_1 = io_now_csr_cycle + 32'h1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 126:37]
  wire [14:0] _T_3 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _funct3_T = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_4 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_5 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:63]
  wire [31:0] _next_reg_T_1 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:63]
  wire [14:0] _T_1084 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_1085 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_48 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_1043 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_1044 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_47 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_1009 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_1010 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_46 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_969 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_970 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_45 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_929 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_930 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_44 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_896 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_897 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_43 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_890 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_891 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_42 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_884 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_885 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_41 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_877 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_878 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_40 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_870 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_871 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_39 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_864 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_865 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_38 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_857 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_858 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_37 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_850 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_851 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_36 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_843 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_844 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_35 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_836 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_837 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_34 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_829 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_830 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_33 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_822 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_823 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_32 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_815 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_816 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_31 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_535 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_536 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_30 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_526 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_527 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_29 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_520 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_521 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_28 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_429 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_430 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_27 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_410 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_411 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_26 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_390 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_391 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_25 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_370 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_371 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_24 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_350 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_351 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_23 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_159 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_160 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_22 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_137 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_21 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_129 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_130 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_20 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_122 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_123 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_19 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_115 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_116 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_18 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_108 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_109 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_17 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_101 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_102 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_16 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_94 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_95 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_15 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_87 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_88 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_14 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_80 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_81 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_13 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_73 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_74 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_12 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_66 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_67 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_11 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_60 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_10 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_56 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_9 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_51 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_52 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_8 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_45 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_46 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_7 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_39 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_40 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_6 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_33 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_34 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_5 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_27 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_28 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_4 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_21 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_22 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_3 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_15 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_16 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_2 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_9 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_10 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_1 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_68 = _T_1 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [4:0] _GEN_139 = _T_7 ? inst[11:7] : _GEN_68; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_210 = _T_13 ? inst[11:7] : _GEN_139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_281 = _T_19 ? inst[11:7] : _GEN_210; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_352 = _T_25 ? inst[11:7] : _GEN_281; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_423 = _T_31 ? inst[11:7] : _GEN_352; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_494 = _T_37 ? inst[11:7] : _GEN_423; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_565 = _T_43 ? inst[11:7] : _GEN_494; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_636 = _T_49 ? inst[11:7] : _GEN_565; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_705 = _T_55 ? inst[11:7] : _GEN_636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_774 = _T_59 ? inst[11:7] : _GEN_705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_878 = _T_63 ? inst[11:7] : _GEN_774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_949 = _T_70 ? inst[11:7] : _GEN_878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1020 = _T_77 ? inst[11:7] : _GEN_949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1091 = _T_84 ? inst[11:7] : _GEN_1020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1162 = _T_91 ? inst[11:7] : _GEN_1091; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1233 = _T_98 ? inst[11:7] : _GEN_1162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1304 = _T_105 ? inst[11:7] : _GEN_1233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1375 = _T_112 ? inst[11:7] : _GEN_1304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1446 = _T_119 ? inst[11:7] : _GEN_1375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1517 = _T_126 ? inst[11:7] : _GEN_1446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1625 = _T_133 ? inst[11:7] : _GEN_1517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1738 = _T_157 ? inst[11:7] : _GEN_1625; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2001 = _T_348 ? inst[11:7] : _GEN_1738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2114 = _T_368 ? inst[11:7] : _GEN_2001; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2227 = _T_388 ? inst[11:7] : _GEN_2114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2305 = _T_408 ? inst[11:7] : _GEN_2227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2418 = _T_427 ? inst[11:7] : _GEN_2305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2518 = _T_518 ? inst[11:7] : _GEN_2418; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2536 = _T_524 ? inst[11:7] : _GEN_2518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2547 = _T_533 ? inst[11:7] : _GEN_2536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2588 = _T_542 ? rs1 : _GEN_2547; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 138:24]
  wire [4:0] _GEN_2838 = _T_593 ? rs1 : _GEN_2588; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 173:22]
  wire [4:0] _GEN_2846 = _T_602 ? rs1 : _GEN_2838; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 179:24]
  wire [4:0] _GEN_2976 = _T_629 ? rs1 : _GEN_2846; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 204:22]
  wire [4:0] _GEN_3048 = _T_647 ? rs1 : _GEN_2976; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 209:23]
  wire [4:0] _GEN_3151 = _T_662 ? rs1 : _GEN_3048; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 215:24]
  wire [4:0] _GEN_3190 = _T_674 ? rs1 : _GEN_3151; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 220:28]
  wire [4:0] _GEN_3299 = _T_702 ? rs1 : _GEN_3190; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 230:24]
  wire [4:0] _GEN_3682 = _T_755 ? rs1 : _GEN_3299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 251:23]
  wire [4:0] _GEN_3752 = _T_767 ? rs1 : _GEN_3682; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 252:23]
  wire [4:0] _GEN_4331 = _T_805 ? rs1 : _GEN_3752; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 259:23]
  wire [4:0] _GEN_4369 = _T_812 ? inst[11:7] : _GEN_4331; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4440 = _T_819 ? inst[11:7] : _GEN_4369; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4511 = _T_826 ? inst[11:7] : _GEN_4440; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4582 = _T_833 ? inst[11:7] : _GEN_4511; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4653 = _T_840 ? inst[11:7] : _GEN_4582; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4724 = _T_847 ? inst[11:7] : _GEN_4653; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4795 = _T_854 ? inst[11:7] : _GEN_4724; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4866 = _T_861 ? inst[11:7] : _GEN_4795; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4915 = _T_868 ? inst[11:7] : _GEN_4866; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4936 = _T_875 ? inst[11:7] : _GEN_4915; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4950 = _T_882 ? inst[11:7] : _GEN_4936; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4957 = _T_888 ? inst[11:7] : _GEN_4950; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5100 = _T_894 ? inst[11:7] : _GEN_4957; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5272 = _T_927 ? inst[11:7] : _GEN_5100; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5444 = _T_967 ? inst[11:7] : _GEN_5272; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5632 = _T_1007 ? inst[11:7] : _GEN_5444; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5804 = _T_1041 ? inst[11:7] : _GEN_5632; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5976 = _T_1082 ? inst[11:7] : _GEN_5804; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rd = io_valid ? _GEN_5976 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [4:0] _GEN_6108 = rd; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [31:0] _next_reg_rd = _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:63]
  wire [31:0] _GEN_32 = 5'h0 == rd ? _T_433 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_33 = 5'h1 == rd ? _T_433 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_34 = 5'h2 == rd ? _T_433 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_35 = 5'h3 == rd ? _T_433 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_36 = 5'h4 == rd ? _T_433 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_37 = 5'h5 == rd ? _T_433 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_38 = 5'h6 == rd ? _T_433 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_39 = 5'h7 == rd ? _T_433 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_40 = 5'h8 == rd ? _T_433 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_41 = 5'h9 == rd ? _T_433 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_42 = 5'ha == rd ? _T_433 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_43 = 5'hb == rd ? _T_433 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_44 = 5'hc == rd ? _T_433 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_45 = 5'hd == rd ? _T_433 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_46 = 5'he == rd ? _T_433 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_47 = 5'hf == rd ? _T_433 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_48 = 5'h10 == rd ? _T_433 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_49 = 5'h11 == rd ? _T_433 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_50 = 5'h12 == rd ? _T_433 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_51 = 5'h13 == rd ? _T_433 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_52 = 5'h14 == rd ? _T_433 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_53 = 5'h15 == rd ? _T_433 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_54 = 5'h16 == rd ? _T_433 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_55 = 5'h17 == rd ? _T_433 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_56 = 5'h18 == rd ? _T_433 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_57 = 5'h19 == rd ? _T_433 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_58 = 5'h1a == rd ? _T_433 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_59 = 5'h1b == rd ? _T_433 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_60 = 5'h1c == rd ? _T_433 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_61 = 5'h1d == rd ? _T_433 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_62 = 5'h1e == rd ? _T_433 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_63 = 5'h1f == rd ? _T_433 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [2:0] _GEN_67 = _T_1 ? inst[14:12] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 18:24]
  wire [6:0] _GEN_69 = _T_1 ? inst[6:0] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 16:24]
  wire [31:0] _GEN_71 = _T_1 ? _GEN_32 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_72 = _T_1 ? _GEN_33 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_73 = _T_1 ? _GEN_34 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_74 = _T_1 ? _GEN_35 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_75 = _T_1 ? _GEN_36 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_76 = _T_1 ? _GEN_37 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_77 = _T_1 ? _GEN_38 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_78 = _T_1 ? _GEN_39 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_79 = _T_1 ? _GEN_40 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_80 = _T_1 ? _GEN_41 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_81 = _T_1 ? _GEN_42 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_82 = _T_1 ? _GEN_43 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_83 = _T_1 ? _GEN_44 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_84 = _T_1 ? _GEN_45 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_85 = _T_1 ? _GEN_46 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_86 = _T_1 ? _GEN_47 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_87 = _T_1 ? _GEN_48 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_88 = _T_1 ? _GEN_49 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_89 = _T_1 ? _GEN_50 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_90 = _T_1 ? _GEN_51 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_91 = _T_1 ? _GEN_52 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_92 = _T_1 ? _GEN_53 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_93 = _T_1 ? _GEN_54 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_94 = _T_1 ? _GEN_55 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_95 = _T_1 ? _GEN_56 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_96 = _T_1 ? _GEN_57 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_97 = _T_1 ? _GEN_58 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_98 = _T_1 ? _GEN_59 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_99 = _T_1 ? _GEN_60 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_100 = _T_1 ? _GEN_61 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_101 = _T_1 ? _GEN_62 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_102 = _T_1 ? _GEN_63 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [2:0] _funct3_T_1 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_11 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_0 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_2 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:67]
  wire [31:0] _next_reg_T_3 = io_valid ? _GEN_5978 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:80]
  wire  _next_reg_T_4 = $signed(_T_300) < $signed(_next_reg_T_3); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:74]
  wire  _next_reg_T_5 = $signed(_T_300) < $signed(_next_reg_T_3); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:74]
  wire [31:0] _next_reg_rd_0 = {{31'd0}, $signed(_T_300) < $signed(_next_reg_T_3)}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_103 = 5'h0 == rd ? _next_reg_rd_0 : _GEN_71; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_104 = 5'h1 == rd ? _next_reg_rd_0 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_105 = 5'h2 == rd ? _next_reg_rd_0 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_106 = 5'h3 == rd ? _next_reg_rd_0 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_107 = 5'h4 == rd ? _next_reg_rd_0 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_108 = 5'h5 == rd ? _next_reg_rd_0 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_109 = 5'h6 == rd ? _next_reg_rd_0 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_110 = 5'h7 == rd ? _next_reg_rd_0 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_111 = 5'h8 == rd ? _next_reg_rd_0 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_112 = 5'h9 == rd ? _next_reg_rd_0 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_113 = 5'ha == rd ? _next_reg_rd_0 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_114 = 5'hb == rd ? _next_reg_rd_0 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_115 = 5'hc == rd ? _next_reg_rd_0 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_116 = 5'hd == rd ? _next_reg_rd_0 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_117 = 5'he == rd ? _next_reg_rd_0 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_118 = 5'hf == rd ? _next_reg_rd_0 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_119 = 5'h10 == rd ? _next_reg_rd_0 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_120 = 5'h11 == rd ? _next_reg_rd_0 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_121 = 5'h12 == rd ? _next_reg_rd_0 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_122 = 5'h13 == rd ? _next_reg_rd_0 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_123 = 5'h14 == rd ? _next_reg_rd_0 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_124 = 5'h15 == rd ? _next_reg_rd_0 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_125 = 5'h16 == rd ? _next_reg_rd_0 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_126 = 5'h17 == rd ? _next_reg_rd_0 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_127 = 5'h18 == rd ? _next_reg_rd_0 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_128 = 5'h19 == rd ? _next_reg_rd_0 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_129 = 5'h1a == rd ? _next_reg_rd_0 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_130 = 5'h1b == rd ? _next_reg_rd_0 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_131 = 5'h1c == rd ? _next_reg_rd_0 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_132 = 5'h1d == rd ? _next_reg_rd_0 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_133 = 5'h1e == rd ? _next_reg_rd_0 : _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_134 = 5'h1f == rd ? _next_reg_rd_0 : _GEN_102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [2:0] _GEN_138 = _T_7 ? inst[14:12] : _GEN_67; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_140 = _T_7 ? inst[6:0] : _GEN_69; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_142 = _T_7 ? _GEN_103 : _GEN_71; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_143 = _T_7 ? _GEN_104 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_144 = _T_7 ? _GEN_105 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_145 = _T_7 ? _GEN_106 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_146 = _T_7 ? _GEN_107 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_147 = _T_7 ? _GEN_108 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_148 = _T_7 ? _GEN_109 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_149 = _T_7 ? _GEN_110 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_150 = _T_7 ? _GEN_111 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_151 = _T_7 ? _GEN_112 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_152 = _T_7 ? _GEN_113 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_153 = _T_7 ? _GEN_114 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_154 = _T_7 ? _GEN_115 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_155 = _T_7 ? _GEN_116 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_156 = _T_7 ? _GEN_117 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_157 = _T_7 ? _GEN_118 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_158 = _T_7 ? _GEN_119 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_159 = _T_7 ? _GEN_120 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_160 = _T_7 ? _GEN_121 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_161 = _T_7 ? _GEN_122 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_162 = _T_7 ? _GEN_123 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_163 = _T_7 ? _GEN_124 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_164 = _T_7 ? _GEN_125 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_165 = _T_7 ? _GEN_126 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_166 = _T_7 ? _GEN_127 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_167 = _T_7 ? _GEN_128 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_168 = _T_7 ? _GEN_129 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_169 = _T_7 ? _GEN_130 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_170 = _T_7 ? _GEN_131 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_171 = _T_7 ? _GEN_132 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_172 = _T_7 ? _GEN_133 : _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_173 = _T_7 ? _GEN_134 : _GEN_102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [2:0] _funct3_T_2 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_17 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_1 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _next_reg_T_6 = _GEN_31 < imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:67]
  wire  _next_reg_T_7 = _GEN_31 < imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:67]
  wire [31:0] _next_reg_rd_1 = {{31'd0}, _GEN_31 < imm}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_174 = 5'h0 == rd ? _next_reg_rd_1 : _GEN_142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_175 = 5'h1 == rd ? _next_reg_rd_1 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_176 = 5'h2 == rd ? _next_reg_rd_1 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_177 = 5'h3 == rd ? _next_reg_rd_1 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_178 = 5'h4 == rd ? _next_reg_rd_1 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_179 = 5'h5 == rd ? _next_reg_rd_1 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_180 = 5'h6 == rd ? _next_reg_rd_1 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_181 = 5'h7 == rd ? _next_reg_rd_1 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_182 = 5'h8 == rd ? _next_reg_rd_1 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_183 = 5'h9 == rd ? _next_reg_rd_1 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_184 = 5'ha == rd ? _next_reg_rd_1 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_185 = 5'hb == rd ? _next_reg_rd_1 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_186 = 5'hc == rd ? _next_reg_rd_1 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_187 = 5'hd == rd ? _next_reg_rd_1 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_188 = 5'he == rd ? _next_reg_rd_1 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_189 = 5'hf == rd ? _next_reg_rd_1 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_190 = 5'h10 == rd ? _next_reg_rd_1 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_191 = 5'h11 == rd ? _next_reg_rd_1 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_192 = 5'h12 == rd ? _next_reg_rd_1 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_193 = 5'h13 == rd ? _next_reg_rd_1 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_194 = 5'h14 == rd ? _next_reg_rd_1 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_195 = 5'h15 == rd ? _next_reg_rd_1 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_196 = 5'h16 == rd ? _next_reg_rd_1 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_197 = 5'h17 == rd ? _next_reg_rd_1 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_198 = 5'h18 == rd ? _next_reg_rd_1 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_199 = 5'h19 == rd ? _next_reg_rd_1 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_200 = 5'h1a == rd ? _next_reg_rd_1 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_201 = 5'h1b == rd ? _next_reg_rd_1 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_202 = 5'h1c == rd ? _next_reg_rd_1 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_203 = 5'h1d == rd ? _next_reg_rd_1 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_204 = 5'h1e == rd ? _next_reg_rd_1 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_205 = 5'h1f == rd ? _next_reg_rd_1 : _GEN_173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [2:0] _GEN_209 = _T_13 ? inst[14:12] : _GEN_138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_211 = _T_13 ? inst[6:0] : _GEN_140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_213 = _T_13 ? _GEN_174 : _GEN_142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_214 = _T_13 ? _GEN_175 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_215 = _T_13 ? _GEN_176 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_216 = _T_13 ? _GEN_177 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_217 = _T_13 ? _GEN_178 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_218 = _T_13 ? _GEN_179 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_219 = _T_13 ? _GEN_180 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_220 = _T_13 ? _GEN_181 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_221 = _T_13 ? _GEN_182 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_222 = _T_13 ? _GEN_183 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_223 = _T_13 ? _GEN_184 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_224 = _T_13 ? _GEN_185 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_225 = _T_13 ? _GEN_186 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_226 = _T_13 ? _GEN_187 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_227 = _T_13 ? _GEN_188 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_228 = _T_13 ? _GEN_189 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_229 = _T_13 ? _GEN_190 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_230 = _T_13 ? _GEN_191 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_231 = _T_13 ? _GEN_192 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_232 = _T_13 ? _GEN_193 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_233 = _T_13 ? _GEN_194 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_234 = _T_13 ? _GEN_195 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_235 = _T_13 ? _GEN_196 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_236 = _T_13 ? _GEN_197 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_237 = _T_13 ? _GEN_198 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_238 = _T_13 ? _GEN_199 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_239 = _T_13 ? _GEN_200 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_240 = _T_13 ? _GEN_201 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_241 = _T_13 ? _GEN_202 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_242 = _T_13 ? _GEN_203 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_243 = _T_13 ? _GEN_204 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_244 = _T_13 ? _GEN_205 : _GEN_173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [2:0] _funct3_T_3 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_23 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_2 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_8 = _GEN_31 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:62]
  wire [31:0] _next_reg_rd_2 = _GEN_31 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:62]
  wire [31:0] _GEN_245 = 5'h0 == rd ? _next_reg_T_8 : _GEN_213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_246 = 5'h1 == rd ? _next_reg_T_8 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_247 = 5'h2 == rd ? _next_reg_T_8 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_248 = 5'h3 == rd ? _next_reg_T_8 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_249 = 5'h4 == rd ? _next_reg_T_8 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_250 = 5'h5 == rd ? _next_reg_T_8 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_251 = 5'h6 == rd ? _next_reg_T_8 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_252 = 5'h7 == rd ? _next_reg_T_8 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_253 = 5'h8 == rd ? _next_reg_T_8 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_254 = 5'h9 == rd ? _next_reg_T_8 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_255 = 5'ha == rd ? _next_reg_T_8 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_256 = 5'hb == rd ? _next_reg_T_8 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_257 = 5'hc == rd ? _next_reg_T_8 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_258 = 5'hd == rd ? _next_reg_T_8 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_259 = 5'he == rd ? _next_reg_T_8 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_260 = 5'hf == rd ? _next_reg_T_8 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_261 = 5'h10 == rd ? _next_reg_T_8 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_262 = 5'h11 == rd ? _next_reg_T_8 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_263 = 5'h12 == rd ? _next_reg_T_8 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_264 = 5'h13 == rd ? _next_reg_T_8 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_265 = 5'h14 == rd ? _next_reg_T_8 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_266 = 5'h15 == rd ? _next_reg_T_8 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_267 = 5'h16 == rd ? _next_reg_T_8 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_268 = 5'h17 == rd ? _next_reg_T_8 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_269 = 5'h18 == rd ? _next_reg_T_8 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_270 = 5'h19 == rd ? _next_reg_T_8 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_271 = 5'h1a == rd ? _next_reg_T_8 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_272 = 5'h1b == rd ? _next_reg_T_8 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_273 = 5'h1c == rd ? _next_reg_T_8 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_274 = 5'h1d == rd ? _next_reg_T_8 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_275 = 5'h1e == rd ? _next_reg_T_8 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_276 = 5'h1f == rd ? _next_reg_T_8 : _GEN_244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [2:0] _GEN_280 = _T_19 ? inst[14:12] : _GEN_209; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_282 = _T_19 ? inst[6:0] : _GEN_211; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_284 = _T_19 ? _GEN_245 : _GEN_213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_285 = _T_19 ? _GEN_246 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_286 = _T_19 ? _GEN_247 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_287 = _T_19 ? _GEN_248 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_288 = _T_19 ? _GEN_249 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_289 = _T_19 ? _GEN_250 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_290 = _T_19 ? _GEN_251 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_291 = _T_19 ? _GEN_252 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_292 = _T_19 ? _GEN_253 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_293 = _T_19 ? _GEN_254 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_294 = _T_19 ? _GEN_255 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_295 = _T_19 ? _GEN_256 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_296 = _T_19 ? _GEN_257 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_297 = _T_19 ? _GEN_258 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_298 = _T_19 ? _GEN_259 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_299 = _T_19 ? _GEN_260 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_300 = _T_19 ? _GEN_261 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_301 = _T_19 ? _GEN_262 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_302 = _T_19 ? _GEN_263 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_303 = _T_19 ? _GEN_264 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_304 = _T_19 ? _GEN_265 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_305 = _T_19 ? _GEN_266 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_306 = _T_19 ? _GEN_267 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_307 = _T_19 ? _GEN_268 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_308 = _T_19 ? _GEN_269 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_309 = _T_19 ? _GEN_270 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_310 = _T_19 ? _GEN_271 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_311 = _T_19 ? _GEN_272 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_312 = _T_19 ? _GEN_273 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_313 = _T_19 ? _GEN_274 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_314 = _T_19 ? _GEN_275 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_315 = _T_19 ? _GEN_276 : _GEN_244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [2:0] _funct3_T_4 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_29 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_3 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_9 = _GEN_31 | imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:62]
  wire [31:0] _next_reg_rd_3 = _GEN_31 | imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:62]
  wire [31:0] _GEN_316 = 5'h0 == rd ? _next_reg_T_9 : _GEN_284; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_317 = 5'h1 == rd ? _next_reg_T_9 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_318 = 5'h2 == rd ? _next_reg_T_9 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_319 = 5'h3 == rd ? _next_reg_T_9 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_320 = 5'h4 == rd ? _next_reg_T_9 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_321 = 5'h5 == rd ? _next_reg_T_9 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_322 = 5'h6 == rd ? _next_reg_T_9 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_323 = 5'h7 == rd ? _next_reg_T_9 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_324 = 5'h8 == rd ? _next_reg_T_9 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_325 = 5'h9 == rd ? _next_reg_T_9 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_326 = 5'ha == rd ? _next_reg_T_9 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_327 = 5'hb == rd ? _next_reg_T_9 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_328 = 5'hc == rd ? _next_reg_T_9 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_329 = 5'hd == rd ? _next_reg_T_9 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_330 = 5'he == rd ? _next_reg_T_9 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_331 = 5'hf == rd ? _next_reg_T_9 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_332 = 5'h10 == rd ? _next_reg_T_9 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_333 = 5'h11 == rd ? _next_reg_T_9 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_334 = 5'h12 == rd ? _next_reg_T_9 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_335 = 5'h13 == rd ? _next_reg_T_9 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_336 = 5'h14 == rd ? _next_reg_T_9 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_337 = 5'h15 == rd ? _next_reg_T_9 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_338 = 5'h16 == rd ? _next_reg_T_9 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_339 = 5'h17 == rd ? _next_reg_T_9 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_340 = 5'h18 == rd ? _next_reg_T_9 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_341 = 5'h19 == rd ? _next_reg_T_9 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_342 = 5'h1a == rd ? _next_reg_T_9 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_343 = 5'h1b == rd ? _next_reg_T_9 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_344 = 5'h1c == rd ? _next_reg_T_9 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_345 = 5'h1d == rd ? _next_reg_T_9 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_346 = 5'h1e == rd ? _next_reg_T_9 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_347 = 5'h1f == rd ? _next_reg_T_9 : _GEN_315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [2:0] _GEN_351 = _T_25 ? inst[14:12] : _GEN_280; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_353 = _T_25 ? inst[6:0] : _GEN_282; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_355 = _T_25 ? _GEN_316 : _GEN_284; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_356 = _T_25 ? _GEN_317 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_357 = _T_25 ? _GEN_318 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_358 = _T_25 ? _GEN_319 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_359 = _T_25 ? _GEN_320 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_360 = _T_25 ? _GEN_321 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_361 = _T_25 ? _GEN_322 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_362 = _T_25 ? _GEN_323 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_363 = _T_25 ? _GEN_324 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_364 = _T_25 ? _GEN_325 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_365 = _T_25 ? _GEN_326 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_366 = _T_25 ? _GEN_327 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_367 = _T_25 ? _GEN_328 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_368 = _T_25 ? _GEN_329 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_369 = _T_25 ? _GEN_330 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_370 = _T_25 ? _GEN_331 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_371 = _T_25 ? _GEN_332 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_372 = _T_25 ? _GEN_333 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_373 = _T_25 ? _GEN_334 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_374 = _T_25 ? _GEN_335 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_375 = _T_25 ? _GEN_336 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_376 = _T_25 ? _GEN_337 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_377 = _T_25 ? _GEN_338 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_378 = _T_25 ? _GEN_339 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_379 = _T_25 ? _GEN_340 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_380 = _T_25 ? _GEN_341 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_381 = _T_25 ? _GEN_342 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_382 = _T_25 ? _GEN_343 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_383 = _T_25 ? _GEN_344 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_384 = _T_25 ? _GEN_345 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_385 = _T_25 ? _GEN_346 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_386 = _T_25 ? _GEN_347 : _GEN_315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [2:0] _funct3_T_5 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_35 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_10 = _GEN_31 ^ imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:62]
  wire [31:0] _next_reg_rd_4 = _GEN_31 ^ imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:62]
  wire [31:0] _GEN_387 = 5'h0 == rd ? _next_reg_T_10 : _GEN_355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_388 = 5'h1 == rd ? _next_reg_T_10 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_389 = 5'h2 == rd ? _next_reg_T_10 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_390 = 5'h3 == rd ? _next_reg_T_10 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_391 = 5'h4 == rd ? _next_reg_T_10 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_392 = 5'h5 == rd ? _next_reg_T_10 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_393 = 5'h6 == rd ? _next_reg_T_10 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_394 = 5'h7 == rd ? _next_reg_T_10 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_395 = 5'h8 == rd ? _next_reg_T_10 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_396 = 5'h9 == rd ? _next_reg_T_10 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_397 = 5'ha == rd ? _next_reg_T_10 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_398 = 5'hb == rd ? _next_reg_T_10 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_399 = 5'hc == rd ? _next_reg_T_10 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_400 = 5'hd == rd ? _next_reg_T_10 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_401 = 5'he == rd ? _next_reg_T_10 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_402 = 5'hf == rd ? _next_reg_T_10 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_403 = 5'h10 == rd ? _next_reg_T_10 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_404 = 5'h11 == rd ? _next_reg_T_10 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_405 = 5'h12 == rd ? _next_reg_T_10 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_406 = 5'h13 == rd ? _next_reg_T_10 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_407 = 5'h14 == rd ? _next_reg_T_10 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_408 = 5'h15 == rd ? _next_reg_T_10 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_409 = 5'h16 == rd ? _next_reg_T_10 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_410 = 5'h17 == rd ? _next_reg_T_10 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_411 = 5'h18 == rd ? _next_reg_T_10 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_412 = 5'h19 == rd ? _next_reg_T_10 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_413 = 5'h1a == rd ? _next_reg_T_10 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_414 = 5'h1b == rd ? _next_reg_T_10 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_415 = 5'h1c == rd ? _next_reg_T_10 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_416 = 5'h1d == rd ? _next_reg_T_10 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_417 = 5'h1e == rd ? _next_reg_T_10 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_418 = 5'h1f == rd ? _next_reg_T_10 : _GEN_386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [2:0] _GEN_422 = _T_31 ? inst[14:12] : _GEN_351; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_424 = _T_31 ? inst[6:0] : _GEN_353; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_426 = _T_31 ? _GEN_387 : _GEN_355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_427 = _T_31 ? _GEN_388 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_428 = _T_31 ? _GEN_389 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_429 = _T_31 ? _GEN_390 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_430 = _T_31 ? _GEN_391 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_431 = _T_31 ? _GEN_392 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_432 = _T_31 ? _GEN_393 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_433 = _T_31 ? _GEN_394 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_434 = _T_31 ? _GEN_395 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_435 = _T_31 ? _GEN_396 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_436 = _T_31 ? _GEN_397 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_437 = _T_31 ? _GEN_398 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_438 = _T_31 ? _GEN_399 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_439 = _T_31 ? _GEN_400 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_440 = _T_31 ? _GEN_401 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_441 = _T_31 ? _GEN_402 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_442 = _T_31 ? _GEN_403 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_443 = _T_31 ? _GEN_404 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_444 = _T_31 ? _GEN_405 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_445 = _T_31 ? _GEN_406 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_446 = _T_31 ? _GEN_407 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_447 = _T_31 ? _GEN_408 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_448 = _T_31 ? _GEN_409 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_449 = _T_31 ? _GEN_410 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_450 = _T_31 ? _GEN_411 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_451 = _T_31 ? _GEN_412 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_452 = _T_31 ? _GEN_413 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_453 = _T_31 ? _GEN_414 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_454 = _T_31 ? _GEN_415 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_455 = _T_31 ? _GEN_416 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_456 = _T_31 ? _GEN_417 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_457 = _T_31 ? _GEN_418 : _GEN_386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [2:0] _funct3_T_6 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_41 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _next_reg_T_11 = imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:68]
  wire [31:0] _now_reg_rs1_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [62:0] _GEN_6217 = {{31'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [62:0] _next_reg_T_12 = _GEN_6217 << imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [31:0] _next_reg_rd_5 = _next_reg_T_12[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_458 = 5'h0 == rd ? _next_reg_T_12[31:0] : _GEN_426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_459 = 5'h1 == rd ? _next_reg_T_12[31:0] : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_460 = 5'h2 == rd ? _next_reg_T_12[31:0] : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_461 = 5'h3 == rd ? _next_reg_T_12[31:0] : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_462 = 5'h4 == rd ? _next_reg_T_12[31:0] : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_463 = 5'h5 == rd ? _next_reg_T_12[31:0] : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_464 = 5'h6 == rd ? _next_reg_T_12[31:0] : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_465 = 5'h7 == rd ? _next_reg_T_12[31:0] : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_466 = 5'h8 == rd ? _next_reg_T_12[31:0] : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_467 = 5'h9 == rd ? _next_reg_T_12[31:0] : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_468 = 5'ha == rd ? _next_reg_T_12[31:0] : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_469 = 5'hb == rd ? _next_reg_T_12[31:0] : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_470 = 5'hc == rd ? _next_reg_T_12[31:0] : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_471 = 5'hd == rd ? _next_reg_T_12[31:0] : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_472 = 5'he == rd ? _next_reg_T_12[31:0] : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_473 = 5'hf == rd ? _next_reg_T_12[31:0] : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_474 = 5'h10 == rd ? _next_reg_T_12[31:0] : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_475 = 5'h11 == rd ? _next_reg_T_12[31:0] : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_476 = 5'h12 == rd ? _next_reg_T_12[31:0] : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_477 = 5'h13 == rd ? _next_reg_T_12[31:0] : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_478 = 5'h14 == rd ? _next_reg_T_12[31:0] : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_479 = 5'h15 == rd ? _next_reg_T_12[31:0] : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_480 = 5'h16 == rd ? _next_reg_T_12[31:0] : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_481 = 5'h17 == rd ? _next_reg_T_12[31:0] : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_482 = 5'h18 == rd ? _next_reg_T_12[31:0] : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_483 = 5'h19 == rd ? _next_reg_T_12[31:0] : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_484 = 5'h1a == rd ? _next_reg_T_12[31:0] : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_485 = 5'h1b == rd ? _next_reg_T_12[31:0] : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_486 = 5'h1c == rd ? _next_reg_T_12[31:0] : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_487 = 5'h1d == rd ? _next_reg_T_12[31:0] : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_488 = 5'h1e == rd ? _next_reg_T_12[31:0] : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_489 = 5'h1f == rd ? _next_reg_T_12[31:0] : _GEN_457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [2:0] _GEN_493 = _T_37 ? inst[14:12] : _GEN_422; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_495 = _T_37 ? inst[6:0] : _GEN_424; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_497 = _T_37 ? _GEN_458 : _GEN_426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_498 = _T_37 ? _GEN_459 : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_499 = _T_37 ? _GEN_460 : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_500 = _T_37 ? _GEN_461 : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_501 = _T_37 ? _GEN_462 : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_502 = _T_37 ? _GEN_463 : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_503 = _T_37 ? _GEN_464 : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_504 = _T_37 ? _GEN_465 : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_505 = _T_37 ? _GEN_466 : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_506 = _T_37 ? _GEN_467 : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_507 = _T_37 ? _GEN_468 : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_508 = _T_37 ? _GEN_469 : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_509 = _T_37 ? _GEN_470 : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_510 = _T_37 ? _GEN_471 : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_511 = _T_37 ? _GEN_472 : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_512 = _T_37 ? _GEN_473 : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_513 = _T_37 ? _GEN_474 : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_514 = _T_37 ? _GEN_475 : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_515 = _T_37 ? _GEN_476 : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_516 = _T_37 ? _GEN_477 : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_517 = _T_37 ? _GEN_478 : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_518 = _T_37 ? _GEN_479 : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_519 = _T_37 ? _GEN_480 : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_520 = _T_37 ? _GEN_481 : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_521 = _T_37 ? _GEN_482 : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_522 = _T_37 ? _GEN_483 : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_523 = _T_37 ? _GEN_484 : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_524 = _T_37 ? _GEN_485 : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_525 = _T_37 ? _GEN_486 : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_526 = _T_37 ? _GEN_487 : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_527 = _T_37 ? _GEN_488 : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_528 = _T_37 ? _GEN_489 : _GEN_457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [2:0] _funct3_T_7 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_47 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _next_reg_T_13 = imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:68]
  wire [31:0] _now_reg_rs1_6 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_14 = _GEN_31 >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:62]
  wire [31:0] _next_reg_rd_6 = _GEN_31 >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:62]
  wire [31:0] _GEN_529 = 5'h0 == rd ? _next_reg_T_14 : _GEN_497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_530 = 5'h1 == rd ? _next_reg_T_14 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_531 = 5'h2 == rd ? _next_reg_T_14 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_532 = 5'h3 == rd ? _next_reg_T_14 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_533 = 5'h4 == rd ? _next_reg_T_14 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_534 = 5'h5 == rd ? _next_reg_T_14 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_535 = 5'h6 == rd ? _next_reg_T_14 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_536 = 5'h7 == rd ? _next_reg_T_14 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_537 = 5'h8 == rd ? _next_reg_T_14 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_538 = 5'h9 == rd ? _next_reg_T_14 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_539 = 5'ha == rd ? _next_reg_T_14 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_540 = 5'hb == rd ? _next_reg_T_14 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_541 = 5'hc == rd ? _next_reg_T_14 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_542 = 5'hd == rd ? _next_reg_T_14 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_543 = 5'he == rd ? _next_reg_T_14 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_544 = 5'hf == rd ? _next_reg_T_14 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_545 = 5'h10 == rd ? _next_reg_T_14 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_546 = 5'h11 == rd ? _next_reg_T_14 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_547 = 5'h12 == rd ? _next_reg_T_14 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_548 = 5'h13 == rd ? _next_reg_T_14 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_549 = 5'h14 == rd ? _next_reg_T_14 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_550 = 5'h15 == rd ? _next_reg_T_14 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_551 = 5'h16 == rd ? _next_reg_T_14 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_552 = 5'h17 == rd ? _next_reg_T_14 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_553 = 5'h18 == rd ? _next_reg_T_14 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_554 = 5'h19 == rd ? _next_reg_T_14 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_555 = 5'h1a == rd ? _next_reg_T_14 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_556 = 5'h1b == rd ? _next_reg_T_14 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_557 = 5'h1c == rd ? _next_reg_T_14 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_558 = 5'h1d == rd ? _next_reg_T_14 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_559 = 5'h1e == rd ? _next_reg_T_14 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_560 = 5'h1f == rd ? _next_reg_T_14 : _GEN_528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [2:0] _GEN_564 = _T_43 ? inst[14:12] : _GEN_493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_566 = _T_43 ? inst[6:0] : _GEN_495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_568 = _T_43 ? _GEN_529 : _GEN_497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_569 = _T_43 ? _GEN_530 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_570 = _T_43 ? _GEN_531 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_571 = _T_43 ? _GEN_532 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_572 = _T_43 ? _GEN_533 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_573 = _T_43 ? _GEN_534 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_574 = _T_43 ? _GEN_535 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_575 = _T_43 ? _GEN_536 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_576 = _T_43 ? _GEN_537 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_577 = _T_43 ? _GEN_538 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_578 = _T_43 ? _GEN_539 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_579 = _T_43 ? _GEN_540 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_580 = _T_43 ? _GEN_541 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_581 = _T_43 ? _GEN_542 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_582 = _T_43 ? _GEN_543 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_583 = _T_43 ? _GEN_544 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_584 = _T_43 ? _GEN_545 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_585 = _T_43 ? _GEN_546 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_586 = _T_43 ? _GEN_547 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_587 = _T_43 ? _GEN_548 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_588 = _T_43 ? _GEN_549 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_589 = _T_43 ? _GEN_550 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_590 = _T_43 ? _GEN_551 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_591 = _T_43 ? _GEN_552 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_592 = _T_43 ? _GEN_553 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_593 = _T_43 ? _GEN_554 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_594 = _T_43 ? _GEN_555 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_595 = _T_43 ? _GEN_556 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_596 = _T_43 ? _GEN_557 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_597 = _T_43 ? _GEN_558 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_598 = _T_43 ? _GEN_559 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_599 = _T_43 ? _GEN_560 : _GEN_528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [2:0] _funct3_T_8 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_53 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_7 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_15 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:63]
  wire [4:0] _next_reg_T_16 = imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:76]
  wire [31:0] _next_reg_T_17 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:70]
  wire [31:0] _next_reg_T_18 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:84]
  wire [31:0] _next_reg_rd_7 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:84]
  wire [31:0] _GEN_600 = 5'h0 == rd ? _next_reg_T_18 : _GEN_568; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_601 = 5'h1 == rd ? _next_reg_T_18 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_602 = 5'h2 == rd ? _next_reg_T_18 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_603 = 5'h3 == rd ? _next_reg_T_18 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_604 = 5'h4 == rd ? _next_reg_T_18 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_605 = 5'h5 == rd ? _next_reg_T_18 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_606 = 5'h6 == rd ? _next_reg_T_18 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_607 = 5'h7 == rd ? _next_reg_T_18 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_608 = 5'h8 == rd ? _next_reg_T_18 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_609 = 5'h9 == rd ? _next_reg_T_18 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_610 = 5'ha == rd ? _next_reg_T_18 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_611 = 5'hb == rd ? _next_reg_T_18 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_612 = 5'hc == rd ? _next_reg_T_18 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_613 = 5'hd == rd ? _next_reg_T_18 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_614 = 5'he == rd ? _next_reg_T_18 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_615 = 5'hf == rd ? _next_reg_T_18 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_616 = 5'h10 == rd ? _next_reg_T_18 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_617 = 5'h11 == rd ? _next_reg_T_18 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_618 = 5'h12 == rd ? _next_reg_T_18 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_619 = 5'h13 == rd ? _next_reg_T_18 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_620 = 5'h14 == rd ? _next_reg_T_18 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_621 = 5'h15 == rd ? _next_reg_T_18 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_622 = 5'h16 == rd ? _next_reg_T_18 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_623 = 5'h17 == rd ? _next_reg_T_18 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_624 = 5'h18 == rd ? _next_reg_T_18 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_625 = 5'h19 == rd ? _next_reg_T_18 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_626 = 5'h1a == rd ? _next_reg_T_18 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_627 = 5'h1b == rd ? _next_reg_T_18 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_628 = 5'h1c == rd ? _next_reg_T_18 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_629 = 5'h1d == rd ? _next_reg_T_18 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_630 = 5'h1e == rd ? _next_reg_T_18 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_631 = 5'h1f == rd ? _next_reg_T_18 : _GEN_599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [2:0] _GEN_635 = _T_49 ? inst[14:12] : _GEN_564; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_637 = _T_49 ? inst[6:0] : _GEN_566; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_639 = _T_49 ? _GEN_600 : _GEN_568; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_640 = _T_49 ? _GEN_601 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_641 = _T_49 ? _GEN_602 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_642 = _T_49 ? _GEN_603 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_643 = _T_49 ? _GEN_604 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_644 = _T_49 ? _GEN_605 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_645 = _T_49 ? _GEN_606 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_646 = _T_49 ? _GEN_607 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_647 = _T_49 ? _GEN_608 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_648 = _T_49 ? _GEN_609 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_649 = _T_49 ? _GEN_610 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_650 = _T_49 ? _GEN_611 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_651 = _T_49 ? _GEN_612 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_652 = _T_49 ? _GEN_613 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_653 = _T_49 ? _GEN_614 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_654 = _T_49 ? _GEN_615 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_655 = _T_49 ? _GEN_616 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_656 = _T_49 ? _GEN_617 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_657 = _T_49 ? _GEN_618 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_658 = _T_49 ? _GEN_619 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_659 = _T_49 ? _GEN_620 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_660 = _T_49 ? _GEN_621 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_661 = _T_49 ? _GEN_622 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_662 = _T_49 ? _GEN_623 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_663 = _T_49 ? _GEN_624 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_664 = _T_49 ? _GEN_625 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_665 = _T_49 ? _GEN_626 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_666 = _T_49 ? _GEN_627 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_667 = _T_49 ? _GEN_628 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_668 = _T_49 ? _GEN_629 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_669 = _T_49 ? _GEN_630 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_670 = _T_49 ? _GEN_631 : _GEN_599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [6:0] _T_57 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  imm_signBit_9 = _imm_T_29[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_rd_8 = imm; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [31:0] _GEN_671 = 5'h0 == rd ? imm : _GEN_639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_672 = 5'h1 == rd ? imm : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_673 = 5'h2 == rd ? imm : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_674 = 5'h3 == rd ? imm : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_675 = 5'h4 == rd ? imm : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_676 = 5'h5 == rd ? imm : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_677 = 5'h6 == rd ? imm : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_678 = 5'h7 == rd ? imm : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_679 = 5'h8 == rd ? imm : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_680 = 5'h9 == rd ? imm : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_681 = 5'ha == rd ? imm : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_682 = 5'hb == rd ? imm : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_683 = 5'hc == rd ? imm : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_684 = 5'hd == rd ? imm : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_685 = 5'he == rd ? imm : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_686 = 5'hf == rd ? imm : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_687 = 5'h10 == rd ? imm : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_688 = 5'h11 == rd ? imm : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_689 = 5'h12 == rd ? imm : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_690 = 5'h13 == rd ? imm : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_691 = 5'h14 == rd ? imm : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_692 = 5'h15 == rd ? imm : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_693 = 5'h16 == rd ? imm : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_694 = 5'h17 == rd ? imm : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_695 = 5'h18 == rd ? imm : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_696 = 5'h19 == rd ? imm : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_697 = 5'h1a == rd ? imm : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_698 = 5'h1b == rd ? imm : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_699 = 5'h1c == rd ? imm : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_700 = 5'h1d == rd ? imm : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_701 = 5'h1e == rd ? imm : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_702 = 5'h1f == rd ? imm : _GEN_670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [6:0] _GEN_706 = _T_55 ? inst[6:0] : _GEN_637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_708 = _T_55 ? _GEN_671 : _GEN_639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_709 = _T_55 ? _GEN_672 : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_710 = _T_55 ? _GEN_673 : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_711 = _T_55 ? _GEN_674 : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_712 = _T_55 ? _GEN_675 : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_713 = _T_55 ? _GEN_676 : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_714 = _T_55 ? _GEN_677 : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_715 = _T_55 ? _GEN_678 : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_716 = _T_55 ? _GEN_679 : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_717 = _T_55 ? _GEN_680 : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_718 = _T_55 ? _GEN_681 : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_719 = _T_55 ? _GEN_682 : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_720 = _T_55 ? _GEN_683 : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_721 = _T_55 ? _GEN_684 : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_722 = _T_55 ? _GEN_685 : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_723 = _T_55 ? _GEN_686 : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_724 = _T_55 ? _GEN_687 : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_725 = _T_55 ? _GEN_688 : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_726 = _T_55 ? _GEN_689 : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_727 = _T_55 ? _GEN_690 : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_728 = _T_55 ? _GEN_691 : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_729 = _T_55 ? _GEN_692 : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_730 = _T_55 ? _GEN_693 : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_731 = _T_55 ? _GEN_694 : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_732 = _T_55 ? _GEN_695 : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_733 = _T_55 ? _GEN_696 : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_734 = _T_55 ? _GEN_697 : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_735 = _T_55 ? _GEN_698 : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_736 = _T_55 ? _GEN_699 : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_737 = _T_55 ? _GEN_700 : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_738 = _T_55 ? _GEN_701 : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_739 = _T_55 ? _GEN_702 : _GEN_670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [6:0] _T_61 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  imm_signBit_10 = _imm_T_29[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [32:0] _next_reg_T_19 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:57]
  wire [31:0] _next_reg_T_20 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:57]
  wire [31:0] _next_reg_rd_9 = _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:57]
  wire [31:0] _GEN_740 = 5'h0 == rd ? _T_334 : _GEN_708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_741 = 5'h1 == rd ? _T_334 : _GEN_709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_742 = 5'h2 == rd ? _T_334 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_743 = 5'h3 == rd ? _T_334 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_744 = 5'h4 == rd ? _T_334 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_745 = 5'h5 == rd ? _T_334 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_746 = 5'h6 == rd ? _T_334 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_747 = 5'h7 == rd ? _T_334 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_748 = 5'h8 == rd ? _T_334 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_749 = 5'h9 == rd ? _T_334 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_750 = 5'ha == rd ? _T_334 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_751 = 5'hb == rd ? _T_334 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_752 = 5'hc == rd ? _T_334 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_753 = 5'hd == rd ? _T_334 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_754 = 5'he == rd ? _T_334 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_755 = 5'hf == rd ? _T_334 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_756 = 5'h10 == rd ? _T_334 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_757 = 5'h11 == rd ? _T_334 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_758 = 5'h12 == rd ? _T_334 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_759 = 5'h13 == rd ? _T_334 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_760 = 5'h14 == rd ? _T_334 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_761 = 5'h15 == rd ? _T_334 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_762 = 5'h16 == rd ? _T_334 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_763 = 5'h17 == rd ? _T_334 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_764 = 5'h18 == rd ? _T_334 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_765 = 5'h19 == rd ? _T_334 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_766 = 5'h1a == rd ? _T_334 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_767 = 5'h1b == rd ? _T_334 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_768 = 5'h1c == rd ? _T_334 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_769 = 5'h1d == rd ? _T_334 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_770 = 5'h1e == rd ? _T_334 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_771 = 5'h1f == rd ? _T_334 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [6:0] _GEN_775 = _T_59 ? inst[6:0] : _GEN_706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_777 = _T_59 ? _GEN_740 : _GEN_708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_778 = _T_59 ? _GEN_741 : _GEN_709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_779 = _T_59 ? _GEN_742 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_780 = _T_59 ? _GEN_743 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_781 = _T_59 ? _GEN_744 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_782 = _T_59 ? _GEN_745 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_783 = _T_59 ? _GEN_746 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_784 = _T_59 ? _GEN_747 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_785 = _T_59 ? _GEN_748 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_786 = _T_59 ? _GEN_749 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_787 = _T_59 ? _GEN_750 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_788 = _T_59 ? _GEN_751 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_789 = _T_59 ? _GEN_752 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_790 = _T_59 ? _GEN_753 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_791 = _T_59 ? _GEN_754 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_792 = _T_59 ? _GEN_755 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_793 = _T_59 ? _GEN_756 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_794 = _T_59 ? _GEN_757 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_795 = _T_59 ? _GEN_758 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_796 = _T_59 ? _GEN_759 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_797 = _T_59 ? _GEN_760 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_798 = _T_59 ? _GEN_761 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_799 = _T_59 ? _GEN_762 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_800 = _T_59 ? _GEN_763 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_801 = _T_59 ? _GEN_764 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_802 = _T_59 ? _GEN_765 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_803 = _T_59 ? _GEN_766 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_804 = _T_59 ? _GEN_767 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_805 = _T_59 ? _GEN_768 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_806 = _T_59 ? _GEN_769 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_807 = _T_59 ? _GEN_770 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_808 = _T_59 ? _GEN_771 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [6:0] _funct7_T = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_9 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_68 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_8 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_21 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [31:0] _next_reg_T_22 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [31:0] _next_reg_rd_10 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [31:0] _GEN_841 = 5'h0 == rd ? _next_reg_T_22 : _GEN_777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_842 = 5'h1 == rd ? _next_reg_T_22 : _GEN_778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_843 = 5'h2 == rd ? _next_reg_T_22 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_844 = 5'h3 == rd ? _next_reg_T_22 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_845 = 5'h4 == rd ? _next_reg_T_22 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_846 = 5'h5 == rd ? _next_reg_T_22 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_847 = 5'h6 == rd ? _next_reg_T_22 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_848 = 5'h7 == rd ? _next_reg_T_22 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_849 = 5'h8 == rd ? _next_reg_T_22 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_850 = 5'h9 == rd ? _next_reg_T_22 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_851 = 5'ha == rd ? _next_reg_T_22 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_852 = 5'hb == rd ? _next_reg_T_22 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_853 = 5'hc == rd ? _next_reg_T_22 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_854 = 5'hd == rd ? _next_reg_T_22 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_855 = 5'he == rd ? _next_reg_T_22 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_856 = 5'hf == rd ? _next_reg_T_22 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_857 = 5'h10 == rd ? _next_reg_T_22 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_858 = 5'h11 == rd ? _next_reg_T_22 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_859 = 5'h12 == rd ? _next_reg_T_22 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_860 = 5'h13 == rd ? _next_reg_T_22 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_861 = 5'h14 == rd ? _next_reg_T_22 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_862 = 5'h15 == rd ? _next_reg_T_22 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_863 = 5'h16 == rd ? _next_reg_T_22 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_864 = 5'h17 == rd ? _next_reg_T_22 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_865 = 5'h18 == rd ? _next_reg_T_22 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_866 = 5'h19 == rd ? _next_reg_T_22 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_867 = 5'h1a == rd ? _next_reg_T_22 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_868 = 5'h1b == rd ? _next_reg_T_22 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_869 = 5'h1c == rd ? _next_reg_T_22 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_870 = 5'h1d == rd ? _next_reg_T_22 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_871 = 5'h1e == rd ? _next_reg_T_22 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_872 = 5'h1f == rd ? _next_reg_T_22 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [6:0] _GEN_874 = _T_63 ? inst[31:25] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 21:24]
  wire [2:0] _GEN_877 = _T_63 ? inst[14:12] : _GEN_635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_879 = _T_63 ? inst[6:0] : _GEN_775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_880 = _T_63 ? _GEN_841 : _GEN_777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_881 = _T_63 ? _GEN_842 : _GEN_778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_882 = _T_63 ? _GEN_843 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_883 = _T_63 ? _GEN_844 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_884 = _T_63 ? _GEN_845 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_885 = _T_63 ? _GEN_846 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_886 = _T_63 ? _GEN_847 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_887 = _T_63 ? _GEN_848 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_888 = _T_63 ? _GEN_849 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_889 = _T_63 ? _GEN_850 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_890 = _T_63 ? _GEN_851 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_891 = _T_63 ? _GEN_852 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_892 = _T_63 ? _GEN_853 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_893 = _T_63 ? _GEN_854 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_894 = _T_63 ? _GEN_855 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_895 = _T_63 ? _GEN_856 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_896 = _T_63 ? _GEN_857 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_897 = _T_63 ? _GEN_858 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_898 = _T_63 ? _GEN_859 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_899 = _T_63 ? _GEN_860 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_900 = _T_63 ? _GEN_861 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_901 = _T_63 ? _GEN_862 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_902 = _T_63 ? _GEN_863 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_903 = _T_63 ? _GEN_864 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_904 = _T_63 ? _GEN_865 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_905 = _T_63 ? _GEN_866 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_906 = _T_63 ? _GEN_867 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_907 = _T_63 ? _GEN_868 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_908 = _T_63 ? _GEN_869 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_909 = _T_63 ? _GEN_870 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_910 = _T_63 ? _GEN_871 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_911 = _T_63 ? _GEN_872 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [6:0] _funct7_T_1 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_10 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_75 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_9 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_23 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:66]
  wire [31:0] _now_reg_rs2_0 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_24 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:88]
  wire  _next_reg_T_25 = $signed(_T_300) < $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:73]
  wire  _next_reg_T_26 = _T_246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:73]
  wire [31:0] _next_reg_rd_11 = {{31'd0}, _T_246}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_912 = 5'h0 == rd ? _next_reg_rd_11 : _GEN_880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_913 = 5'h1 == rd ? _next_reg_rd_11 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_914 = 5'h2 == rd ? _next_reg_rd_11 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_915 = 5'h3 == rd ? _next_reg_rd_11 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_916 = 5'h4 == rd ? _next_reg_rd_11 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_917 = 5'h5 == rd ? _next_reg_rd_11 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_918 = 5'h6 == rd ? _next_reg_rd_11 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_919 = 5'h7 == rd ? _next_reg_rd_11 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_920 = 5'h8 == rd ? _next_reg_rd_11 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_921 = 5'h9 == rd ? _next_reg_rd_11 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_922 = 5'ha == rd ? _next_reg_rd_11 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_923 = 5'hb == rd ? _next_reg_rd_11 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_924 = 5'hc == rd ? _next_reg_rd_11 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_925 = 5'hd == rd ? _next_reg_rd_11 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_926 = 5'he == rd ? _next_reg_rd_11 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_927 = 5'hf == rd ? _next_reg_rd_11 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_928 = 5'h10 == rd ? _next_reg_rd_11 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_929 = 5'h11 == rd ? _next_reg_rd_11 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_930 = 5'h12 == rd ? _next_reg_rd_11 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_931 = 5'h13 == rd ? _next_reg_rd_11 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_932 = 5'h14 == rd ? _next_reg_rd_11 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_933 = 5'h15 == rd ? _next_reg_rd_11 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_934 = 5'h16 == rd ? _next_reg_rd_11 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_935 = 5'h17 == rd ? _next_reg_rd_11 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_936 = 5'h18 == rd ? _next_reg_rd_11 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_937 = 5'h19 == rd ? _next_reg_rd_11 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_938 = 5'h1a == rd ? _next_reg_rd_11 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_939 = 5'h1b == rd ? _next_reg_rd_11 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_940 = 5'h1c == rd ? _next_reg_rd_11 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_941 = 5'h1d == rd ? _next_reg_rd_11 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_942 = 5'h1e == rd ? _next_reg_rd_11 : _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_943 = 5'h1f == rd ? _next_reg_rd_11 : _GEN_911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [6:0] _GEN_945 = _T_70 ? inst[31:25] : _GEN_874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_948 = _T_70 ? inst[14:12] : _GEN_877; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_950 = _T_70 ? inst[6:0] : _GEN_879; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_951 = _T_70 ? _GEN_912 : _GEN_880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_952 = _T_70 ? _GEN_913 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_953 = _T_70 ? _GEN_914 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_954 = _T_70 ? _GEN_915 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_955 = _T_70 ? _GEN_916 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_956 = _T_70 ? _GEN_917 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_957 = _T_70 ? _GEN_918 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_958 = _T_70 ? _GEN_919 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_959 = _T_70 ? _GEN_920 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_960 = _T_70 ? _GEN_921 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_961 = _T_70 ? _GEN_922 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_962 = _T_70 ? _GEN_923 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_963 = _T_70 ? _GEN_924 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_964 = _T_70 ? _GEN_925 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_965 = _T_70 ? _GEN_926 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_966 = _T_70 ? _GEN_927 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_967 = _T_70 ? _GEN_928 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_968 = _T_70 ? _GEN_929 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_969 = _T_70 ? _GEN_930 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_970 = _T_70 ? _GEN_931 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_971 = _T_70 ? _GEN_932 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_972 = _T_70 ? _GEN_933 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_973 = _T_70 ? _GEN_934 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_974 = _T_70 ? _GEN_935 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_975 = _T_70 ? _GEN_936 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_976 = _T_70 ? _GEN_937 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_977 = _T_70 ? _GEN_938 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_978 = _T_70 ? _GEN_939 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_979 = _T_70 ? _GEN_940 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_980 = _T_70 ? _GEN_941 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_981 = _T_70 ? _GEN_942 : _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_982 = _T_70 ? _GEN_943 : _GEN_911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [6:0] _funct7_T_2 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_11 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_82 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_10 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_1 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_27 = _GEN_31 < _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:66]
  wire  _next_reg_T_28 = _T_273; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:66]
  wire [31:0] _next_reg_rd_12 = {{31'd0}, _T_273}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_983 = 5'h0 == rd ? _next_reg_rd_12 : _GEN_951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_984 = 5'h1 == rd ? _next_reg_rd_12 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_985 = 5'h2 == rd ? _next_reg_rd_12 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_986 = 5'h3 == rd ? _next_reg_rd_12 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_987 = 5'h4 == rd ? _next_reg_rd_12 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_988 = 5'h5 == rd ? _next_reg_rd_12 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_989 = 5'h6 == rd ? _next_reg_rd_12 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_990 = 5'h7 == rd ? _next_reg_rd_12 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_991 = 5'h8 == rd ? _next_reg_rd_12 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_992 = 5'h9 == rd ? _next_reg_rd_12 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_993 = 5'ha == rd ? _next_reg_rd_12 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_994 = 5'hb == rd ? _next_reg_rd_12 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_995 = 5'hc == rd ? _next_reg_rd_12 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_996 = 5'hd == rd ? _next_reg_rd_12 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_997 = 5'he == rd ? _next_reg_rd_12 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_998 = 5'hf == rd ? _next_reg_rd_12 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_999 = 5'h10 == rd ? _next_reg_rd_12 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1000 = 5'h11 == rd ? _next_reg_rd_12 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1001 = 5'h12 == rd ? _next_reg_rd_12 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1002 = 5'h13 == rd ? _next_reg_rd_12 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1003 = 5'h14 == rd ? _next_reg_rd_12 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1004 = 5'h15 == rd ? _next_reg_rd_12 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1005 = 5'h16 == rd ? _next_reg_rd_12 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1006 = 5'h17 == rd ? _next_reg_rd_12 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1007 = 5'h18 == rd ? _next_reg_rd_12 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1008 = 5'h19 == rd ? _next_reg_rd_12 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1009 = 5'h1a == rd ? _next_reg_rd_12 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1010 = 5'h1b == rd ? _next_reg_rd_12 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1011 = 5'h1c == rd ? _next_reg_rd_12 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1012 = 5'h1d == rd ? _next_reg_rd_12 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1013 = 5'h1e == rd ? _next_reg_rd_12 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1014 = 5'h1f == rd ? _next_reg_rd_12 : _GEN_982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [6:0] _GEN_1016 = _T_77 ? inst[31:25] : _GEN_945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1019 = _T_77 ? inst[14:12] : _GEN_948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1021 = _T_77 ? inst[6:0] : _GEN_950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1022 = _T_77 ? _GEN_983 : _GEN_951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1023 = _T_77 ? _GEN_984 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1024 = _T_77 ? _GEN_985 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1025 = _T_77 ? _GEN_986 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1026 = _T_77 ? _GEN_987 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1027 = _T_77 ? _GEN_988 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1028 = _T_77 ? _GEN_989 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1029 = _T_77 ? _GEN_990 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1030 = _T_77 ? _GEN_991 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1031 = _T_77 ? _GEN_992 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1032 = _T_77 ? _GEN_993 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1033 = _T_77 ? _GEN_994 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1034 = _T_77 ? _GEN_995 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1035 = _T_77 ? _GEN_996 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1036 = _T_77 ? _GEN_997 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1037 = _T_77 ? _GEN_998 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1038 = _T_77 ? _GEN_999 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1039 = _T_77 ? _GEN_1000 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1040 = _T_77 ? _GEN_1001 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1041 = _T_77 ? _GEN_1002 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1042 = _T_77 ? _GEN_1003 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1043 = _T_77 ? _GEN_1004 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1044 = _T_77 ? _GEN_1005 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1045 = _T_77 ? _GEN_1006 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1046 = _T_77 ? _GEN_1007 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1047 = _T_77 ? _GEN_1008 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1048 = _T_77 ? _GEN_1009 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1049 = _T_77 ? _GEN_1010 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1050 = _T_77 ? _GEN_1011 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1051 = _T_77 ? _GEN_1012 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1052 = _T_77 ? _GEN_1013 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1053 = _T_77 ? _GEN_1014 : _GEN_982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [6:0] _funct7_T_3 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_12 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_89 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_11 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_2 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_29 = _GEN_31 & _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:61]
  wire [31:0] _next_reg_rd_13 = _GEN_31 & _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:61]
  wire [31:0] _GEN_1054 = 5'h0 == rd ? _next_reg_T_29 : _GEN_1022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1055 = 5'h1 == rd ? _next_reg_T_29 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1056 = 5'h2 == rd ? _next_reg_T_29 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1057 = 5'h3 == rd ? _next_reg_T_29 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1058 = 5'h4 == rd ? _next_reg_T_29 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1059 = 5'h5 == rd ? _next_reg_T_29 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1060 = 5'h6 == rd ? _next_reg_T_29 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1061 = 5'h7 == rd ? _next_reg_T_29 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1062 = 5'h8 == rd ? _next_reg_T_29 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1063 = 5'h9 == rd ? _next_reg_T_29 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1064 = 5'ha == rd ? _next_reg_T_29 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1065 = 5'hb == rd ? _next_reg_T_29 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1066 = 5'hc == rd ? _next_reg_T_29 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1067 = 5'hd == rd ? _next_reg_T_29 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1068 = 5'he == rd ? _next_reg_T_29 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1069 = 5'hf == rd ? _next_reg_T_29 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1070 = 5'h10 == rd ? _next_reg_T_29 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1071 = 5'h11 == rd ? _next_reg_T_29 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1072 = 5'h12 == rd ? _next_reg_T_29 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1073 = 5'h13 == rd ? _next_reg_T_29 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1074 = 5'h14 == rd ? _next_reg_T_29 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1075 = 5'h15 == rd ? _next_reg_T_29 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1076 = 5'h16 == rd ? _next_reg_T_29 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1077 = 5'h17 == rd ? _next_reg_T_29 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1078 = 5'h18 == rd ? _next_reg_T_29 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1079 = 5'h19 == rd ? _next_reg_T_29 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1080 = 5'h1a == rd ? _next_reg_T_29 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1081 = 5'h1b == rd ? _next_reg_T_29 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1082 = 5'h1c == rd ? _next_reg_T_29 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1083 = 5'h1d == rd ? _next_reg_T_29 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1084 = 5'h1e == rd ? _next_reg_T_29 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1085 = 5'h1f == rd ? _next_reg_T_29 : _GEN_1053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [6:0] _GEN_1087 = _T_84 ? inst[31:25] : _GEN_1016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1090 = _T_84 ? inst[14:12] : _GEN_1019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1092 = _T_84 ? inst[6:0] : _GEN_1021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1093 = _T_84 ? _GEN_1054 : _GEN_1022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1094 = _T_84 ? _GEN_1055 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1095 = _T_84 ? _GEN_1056 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1096 = _T_84 ? _GEN_1057 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1097 = _T_84 ? _GEN_1058 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1098 = _T_84 ? _GEN_1059 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1099 = _T_84 ? _GEN_1060 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1100 = _T_84 ? _GEN_1061 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1101 = _T_84 ? _GEN_1062 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1102 = _T_84 ? _GEN_1063 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1103 = _T_84 ? _GEN_1064 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1104 = _T_84 ? _GEN_1065 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1105 = _T_84 ? _GEN_1066 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1106 = _T_84 ? _GEN_1067 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1107 = _T_84 ? _GEN_1068 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1108 = _T_84 ? _GEN_1069 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1109 = _T_84 ? _GEN_1070 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1110 = _T_84 ? _GEN_1071 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1111 = _T_84 ? _GEN_1072 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1112 = _T_84 ? _GEN_1073 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1113 = _T_84 ? _GEN_1074 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1114 = _T_84 ? _GEN_1075 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1115 = _T_84 ? _GEN_1076 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1116 = _T_84 ? _GEN_1077 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1117 = _T_84 ? _GEN_1078 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1118 = _T_84 ? _GEN_1079 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1119 = _T_84 ? _GEN_1080 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1120 = _T_84 ? _GEN_1081 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1121 = _T_84 ? _GEN_1082 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1122 = _T_84 ? _GEN_1083 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1123 = _T_84 ? _GEN_1084 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1124 = _T_84 ? _GEN_1085 : _GEN_1053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [6:0] _funct7_T_4 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_13 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_96 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_12 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_3 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_30 = _GEN_31 | _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:61]
  wire [31:0] _next_reg_rd_14 = _GEN_31 | _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:61]
  wire [31:0] _GEN_1125 = 5'h0 == rd ? _next_reg_T_30 : _GEN_1093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1126 = 5'h1 == rd ? _next_reg_T_30 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1127 = 5'h2 == rd ? _next_reg_T_30 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1128 = 5'h3 == rd ? _next_reg_T_30 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1129 = 5'h4 == rd ? _next_reg_T_30 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1130 = 5'h5 == rd ? _next_reg_T_30 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1131 = 5'h6 == rd ? _next_reg_T_30 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1132 = 5'h7 == rd ? _next_reg_T_30 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1133 = 5'h8 == rd ? _next_reg_T_30 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1134 = 5'h9 == rd ? _next_reg_T_30 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1135 = 5'ha == rd ? _next_reg_T_30 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1136 = 5'hb == rd ? _next_reg_T_30 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1137 = 5'hc == rd ? _next_reg_T_30 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1138 = 5'hd == rd ? _next_reg_T_30 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1139 = 5'he == rd ? _next_reg_T_30 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1140 = 5'hf == rd ? _next_reg_T_30 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1141 = 5'h10 == rd ? _next_reg_T_30 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1142 = 5'h11 == rd ? _next_reg_T_30 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1143 = 5'h12 == rd ? _next_reg_T_30 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1144 = 5'h13 == rd ? _next_reg_T_30 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1145 = 5'h14 == rd ? _next_reg_T_30 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1146 = 5'h15 == rd ? _next_reg_T_30 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1147 = 5'h16 == rd ? _next_reg_T_30 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1148 = 5'h17 == rd ? _next_reg_T_30 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1149 = 5'h18 == rd ? _next_reg_T_30 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1150 = 5'h19 == rd ? _next_reg_T_30 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1151 = 5'h1a == rd ? _next_reg_T_30 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1152 = 5'h1b == rd ? _next_reg_T_30 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1153 = 5'h1c == rd ? _next_reg_T_30 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1154 = 5'h1d == rd ? _next_reg_T_30 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1155 = 5'h1e == rd ? _next_reg_T_30 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1156 = 5'h1f == rd ? _next_reg_T_30 : _GEN_1124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [6:0] _GEN_1158 = _T_91 ? inst[31:25] : _GEN_1087; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1161 = _T_91 ? inst[14:12] : _GEN_1090; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1163 = _T_91 ? inst[6:0] : _GEN_1092; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1164 = _T_91 ? _GEN_1125 : _GEN_1093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1165 = _T_91 ? _GEN_1126 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1166 = _T_91 ? _GEN_1127 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1167 = _T_91 ? _GEN_1128 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1168 = _T_91 ? _GEN_1129 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1169 = _T_91 ? _GEN_1130 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1170 = _T_91 ? _GEN_1131 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1171 = _T_91 ? _GEN_1132 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1172 = _T_91 ? _GEN_1133 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1173 = _T_91 ? _GEN_1134 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1174 = _T_91 ? _GEN_1135 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1175 = _T_91 ? _GEN_1136 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1176 = _T_91 ? _GEN_1137 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1177 = _T_91 ? _GEN_1138 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1178 = _T_91 ? _GEN_1139 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1179 = _T_91 ? _GEN_1140 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1180 = _T_91 ? _GEN_1141 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1181 = _T_91 ? _GEN_1142 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1182 = _T_91 ? _GEN_1143 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1183 = _T_91 ? _GEN_1144 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1184 = _T_91 ? _GEN_1145 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1185 = _T_91 ? _GEN_1146 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1186 = _T_91 ? _GEN_1147 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1187 = _T_91 ? _GEN_1148 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1188 = _T_91 ? _GEN_1149 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1189 = _T_91 ? _GEN_1150 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1190 = _T_91 ? _GEN_1151 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1191 = _T_91 ? _GEN_1152 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1192 = _T_91 ? _GEN_1153 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1193 = _T_91 ? _GEN_1154 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1194 = _T_91 ? _GEN_1155 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1195 = _T_91 ? _GEN_1156 : _GEN_1124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [6:0] _funct7_T_5 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_14 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_103 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_13 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_4 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_31 = _GEN_31 ^ _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:61]
  wire [31:0] _next_reg_rd_15 = _GEN_31 ^ _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:61]
  wire [31:0] _GEN_1196 = 5'h0 == rd ? _next_reg_T_31 : _GEN_1164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1197 = 5'h1 == rd ? _next_reg_T_31 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1198 = 5'h2 == rd ? _next_reg_T_31 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1199 = 5'h3 == rd ? _next_reg_T_31 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1200 = 5'h4 == rd ? _next_reg_T_31 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1201 = 5'h5 == rd ? _next_reg_T_31 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1202 = 5'h6 == rd ? _next_reg_T_31 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1203 = 5'h7 == rd ? _next_reg_T_31 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1204 = 5'h8 == rd ? _next_reg_T_31 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1205 = 5'h9 == rd ? _next_reg_T_31 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1206 = 5'ha == rd ? _next_reg_T_31 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1207 = 5'hb == rd ? _next_reg_T_31 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1208 = 5'hc == rd ? _next_reg_T_31 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1209 = 5'hd == rd ? _next_reg_T_31 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1210 = 5'he == rd ? _next_reg_T_31 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1211 = 5'hf == rd ? _next_reg_T_31 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1212 = 5'h10 == rd ? _next_reg_T_31 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1213 = 5'h11 == rd ? _next_reg_T_31 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1214 = 5'h12 == rd ? _next_reg_T_31 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1215 = 5'h13 == rd ? _next_reg_T_31 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1216 = 5'h14 == rd ? _next_reg_T_31 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1217 = 5'h15 == rd ? _next_reg_T_31 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1218 = 5'h16 == rd ? _next_reg_T_31 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1219 = 5'h17 == rd ? _next_reg_T_31 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1220 = 5'h18 == rd ? _next_reg_T_31 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1221 = 5'h19 == rd ? _next_reg_T_31 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1222 = 5'h1a == rd ? _next_reg_T_31 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1223 = 5'h1b == rd ? _next_reg_T_31 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1224 = 5'h1c == rd ? _next_reg_T_31 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1225 = 5'h1d == rd ? _next_reg_T_31 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1226 = 5'h1e == rd ? _next_reg_T_31 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1227 = 5'h1f == rd ? _next_reg_T_31 : _GEN_1195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [6:0] _GEN_1229 = _T_98 ? inst[31:25] : _GEN_1158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1232 = _T_98 ? inst[14:12] : _GEN_1161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1234 = _T_98 ? inst[6:0] : _GEN_1163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1235 = _T_98 ? _GEN_1196 : _GEN_1164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1236 = _T_98 ? _GEN_1197 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1237 = _T_98 ? _GEN_1198 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1238 = _T_98 ? _GEN_1199 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1239 = _T_98 ? _GEN_1200 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1240 = _T_98 ? _GEN_1201 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1241 = _T_98 ? _GEN_1202 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1242 = _T_98 ? _GEN_1203 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1243 = _T_98 ? _GEN_1204 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1244 = _T_98 ? _GEN_1205 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1245 = _T_98 ? _GEN_1206 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1246 = _T_98 ? _GEN_1207 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1247 = _T_98 ? _GEN_1208 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1248 = _T_98 ? _GEN_1209 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1249 = _T_98 ? _GEN_1210 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1250 = _T_98 ? _GEN_1211 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1251 = _T_98 ? _GEN_1212 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1252 = _T_98 ? _GEN_1213 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1253 = _T_98 ? _GEN_1214 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1254 = _T_98 ? _GEN_1215 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1255 = _T_98 ? _GEN_1216 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1256 = _T_98 ? _GEN_1217 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1257 = _T_98 ? _GEN_1218 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1258 = _T_98 ? _GEN_1219 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1259 = _T_98 ? _GEN_1220 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1260 = _T_98 ? _GEN_1221 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1261 = _T_98 ? _GEN_1222 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1262 = _T_98 ? _GEN_1223 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1263 = _T_98 ? _GEN_1224 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1264 = _T_98 ? _GEN_1225 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1265 = _T_98 ? _GEN_1226 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1266 = _T_98 ? _GEN_1227 : _GEN_1195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [6:0] _funct7_T_6 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_15 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_110 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs2_5 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [4:0] _next_reg_T_32 = _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:76]
  wire [31:0] _now_reg_rs1_14 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [62:0] _GEN_6218 = {{31'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [62:0] _next_reg_T_33 = _GEN_6218 << _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [31:0] _next_reg_rd_16 = _next_reg_T_33[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1267 = 5'h0 == rd ? _next_reg_T_33[31:0] : _GEN_1235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1268 = 5'h1 == rd ? _next_reg_T_33[31:0] : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1269 = 5'h2 == rd ? _next_reg_T_33[31:0] : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1270 = 5'h3 == rd ? _next_reg_T_33[31:0] : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1271 = 5'h4 == rd ? _next_reg_T_33[31:0] : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1272 = 5'h5 == rd ? _next_reg_T_33[31:0] : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1273 = 5'h6 == rd ? _next_reg_T_33[31:0] : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1274 = 5'h7 == rd ? _next_reg_T_33[31:0] : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1275 = 5'h8 == rd ? _next_reg_T_33[31:0] : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1276 = 5'h9 == rd ? _next_reg_T_33[31:0] : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1277 = 5'ha == rd ? _next_reg_T_33[31:0] : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1278 = 5'hb == rd ? _next_reg_T_33[31:0] : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1279 = 5'hc == rd ? _next_reg_T_33[31:0] : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1280 = 5'hd == rd ? _next_reg_T_33[31:0] : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1281 = 5'he == rd ? _next_reg_T_33[31:0] : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1282 = 5'hf == rd ? _next_reg_T_33[31:0] : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1283 = 5'h10 == rd ? _next_reg_T_33[31:0] : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1284 = 5'h11 == rd ? _next_reg_T_33[31:0] : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1285 = 5'h12 == rd ? _next_reg_T_33[31:0] : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1286 = 5'h13 == rd ? _next_reg_T_33[31:0] : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1287 = 5'h14 == rd ? _next_reg_T_33[31:0] : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1288 = 5'h15 == rd ? _next_reg_T_33[31:0] : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1289 = 5'h16 == rd ? _next_reg_T_33[31:0] : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1290 = 5'h17 == rd ? _next_reg_T_33[31:0] : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1291 = 5'h18 == rd ? _next_reg_T_33[31:0] : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1292 = 5'h19 == rd ? _next_reg_T_33[31:0] : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1293 = 5'h1a == rd ? _next_reg_T_33[31:0] : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1294 = 5'h1b == rd ? _next_reg_T_33[31:0] : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1295 = 5'h1c == rd ? _next_reg_T_33[31:0] : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1296 = 5'h1d == rd ? _next_reg_T_33[31:0] : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1297 = 5'h1e == rd ? _next_reg_T_33[31:0] : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1298 = 5'h1f == rd ? _next_reg_T_33[31:0] : _GEN_1266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [6:0] _GEN_1300 = _T_105 ? inst[31:25] : _GEN_1229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1303 = _T_105 ? inst[14:12] : _GEN_1232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1305 = _T_105 ? inst[6:0] : _GEN_1234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1306 = _T_105 ? _GEN_1267 : _GEN_1235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1307 = _T_105 ? _GEN_1268 : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1308 = _T_105 ? _GEN_1269 : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1309 = _T_105 ? _GEN_1270 : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1310 = _T_105 ? _GEN_1271 : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1311 = _T_105 ? _GEN_1272 : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1312 = _T_105 ? _GEN_1273 : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1313 = _T_105 ? _GEN_1274 : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1314 = _T_105 ? _GEN_1275 : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1315 = _T_105 ? _GEN_1276 : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1316 = _T_105 ? _GEN_1277 : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1317 = _T_105 ? _GEN_1278 : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1318 = _T_105 ? _GEN_1279 : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1319 = _T_105 ? _GEN_1280 : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1320 = _T_105 ? _GEN_1281 : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1321 = _T_105 ? _GEN_1282 : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1322 = _T_105 ? _GEN_1283 : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1323 = _T_105 ? _GEN_1284 : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1324 = _T_105 ? _GEN_1285 : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1325 = _T_105 ? _GEN_1286 : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1326 = _T_105 ? _GEN_1287 : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1327 = _T_105 ? _GEN_1288 : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1328 = _T_105 ? _GEN_1289 : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1329 = _T_105 ? _GEN_1290 : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1330 = _T_105 ? _GEN_1291 : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1331 = _T_105 ? _GEN_1292 : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1332 = _T_105 ? _GEN_1293 : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1333 = _T_105 ? _GEN_1294 : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1334 = _T_105 ? _GEN_1295 : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1335 = _T_105 ? _GEN_1296 : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1336 = _T_105 ? _GEN_1297 : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1337 = _T_105 ? _GEN_1298 : _GEN_1266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [6:0] _funct7_T_7 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_16 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_117 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs2_6 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [4:0] _next_reg_T_34 = _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:76]
  wire [31:0] _now_reg_rs1_15 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_35 = _GEN_31 >> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:61]
  wire [31:0] _next_reg_rd_17 = _GEN_31 >> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:61]
  wire [31:0] _GEN_1338 = 5'h0 == rd ? _next_reg_T_35 : _GEN_1306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1339 = 5'h1 == rd ? _next_reg_T_35 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1340 = 5'h2 == rd ? _next_reg_T_35 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1341 = 5'h3 == rd ? _next_reg_T_35 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1342 = 5'h4 == rd ? _next_reg_T_35 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1343 = 5'h5 == rd ? _next_reg_T_35 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1344 = 5'h6 == rd ? _next_reg_T_35 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1345 = 5'h7 == rd ? _next_reg_T_35 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1346 = 5'h8 == rd ? _next_reg_T_35 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1347 = 5'h9 == rd ? _next_reg_T_35 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1348 = 5'ha == rd ? _next_reg_T_35 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1349 = 5'hb == rd ? _next_reg_T_35 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1350 = 5'hc == rd ? _next_reg_T_35 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1351 = 5'hd == rd ? _next_reg_T_35 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1352 = 5'he == rd ? _next_reg_T_35 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1353 = 5'hf == rd ? _next_reg_T_35 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1354 = 5'h10 == rd ? _next_reg_T_35 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1355 = 5'h11 == rd ? _next_reg_T_35 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1356 = 5'h12 == rd ? _next_reg_T_35 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1357 = 5'h13 == rd ? _next_reg_T_35 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1358 = 5'h14 == rd ? _next_reg_T_35 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1359 = 5'h15 == rd ? _next_reg_T_35 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1360 = 5'h16 == rd ? _next_reg_T_35 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1361 = 5'h17 == rd ? _next_reg_T_35 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1362 = 5'h18 == rd ? _next_reg_T_35 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1363 = 5'h19 == rd ? _next_reg_T_35 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1364 = 5'h1a == rd ? _next_reg_T_35 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1365 = 5'h1b == rd ? _next_reg_T_35 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1366 = 5'h1c == rd ? _next_reg_T_35 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1367 = 5'h1d == rd ? _next_reg_T_35 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1368 = 5'h1e == rd ? _next_reg_T_35 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1369 = 5'h1f == rd ? _next_reg_T_35 : _GEN_1337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [6:0] _GEN_1371 = _T_112 ? inst[31:25] : _GEN_1300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1374 = _T_112 ? inst[14:12] : _GEN_1303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1376 = _T_112 ? inst[6:0] : _GEN_1305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1377 = _T_112 ? _GEN_1338 : _GEN_1306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1378 = _T_112 ? _GEN_1339 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1379 = _T_112 ? _GEN_1340 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1380 = _T_112 ? _GEN_1341 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1381 = _T_112 ? _GEN_1342 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1382 = _T_112 ? _GEN_1343 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1383 = _T_112 ? _GEN_1344 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1384 = _T_112 ? _GEN_1345 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1385 = _T_112 ? _GEN_1346 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1386 = _T_112 ? _GEN_1347 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1387 = _T_112 ? _GEN_1348 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1388 = _T_112 ? _GEN_1349 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1389 = _T_112 ? _GEN_1350 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1390 = _T_112 ? _GEN_1351 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1391 = _T_112 ? _GEN_1352 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1392 = _T_112 ? _GEN_1353 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1393 = _T_112 ? _GEN_1354 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1394 = _T_112 ? _GEN_1355 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1395 = _T_112 ? _GEN_1356 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1396 = _T_112 ? _GEN_1357 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1397 = _T_112 ? _GEN_1358 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1398 = _T_112 ? _GEN_1359 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1399 = _T_112 ? _GEN_1360 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1400 = _T_112 ? _GEN_1361 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1401 = _T_112 ? _GEN_1362 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1402 = _T_112 ? _GEN_1363 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1403 = _T_112 ? _GEN_1364 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1404 = _T_112 ? _GEN_1365 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1405 = _T_112 ? _GEN_1366 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1406 = _T_112 ? _GEN_1367 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1407 = _T_112 ? _GEN_1368 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1408 = _T_112 ? _GEN_1369 : _GEN_1337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [6:0] _funct7_T_8 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_17 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_124 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_16 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_7 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_36 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [31:0] _next_reg_T_37 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [31:0] _next_reg_rd_18 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [31:0] _GEN_1409 = 5'h0 == rd ? _next_reg_T_37 : _GEN_1377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1410 = 5'h1 == rd ? _next_reg_T_37 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1411 = 5'h2 == rd ? _next_reg_T_37 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1412 = 5'h3 == rd ? _next_reg_T_37 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1413 = 5'h4 == rd ? _next_reg_T_37 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1414 = 5'h5 == rd ? _next_reg_T_37 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1415 = 5'h6 == rd ? _next_reg_T_37 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1416 = 5'h7 == rd ? _next_reg_T_37 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1417 = 5'h8 == rd ? _next_reg_T_37 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1418 = 5'h9 == rd ? _next_reg_T_37 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1419 = 5'ha == rd ? _next_reg_T_37 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1420 = 5'hb == rd ? _next_reg_T_37 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1421 = 5'hc == rd ? _next_reg_T_37 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1422 = 5'hd == rd ? _next_reg_T_37 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1423 = 5'he == rd ? _next_reg_T_37 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1424 = 5'hf == rd ? _next_reg_T_37 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1425 = 5'h10 == rd ? _next_reg_T_37 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1426 = 5'h11 == rd ? _next_reg_T_37 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1427 = 5'h12 == rd ? _next_reg_T_37 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1428 = 5'h13 == rd ? _next_reg_T_37 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1429 = 5'h14 == rd ? _next_reg_T_37 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1430 = 5'h15 == rd ? _next_reg_T_37 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1431 = 5'h16 == rd ? _next_reg_T_37 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1432 = 5'h17 == rd ? _next_reg_T_37 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1433 = 5'h18 == rd ? _next_reg_T_37 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1434 = 5'h19 == rd ? _next_reg_T_37 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1435 = 5'h1a == rd ? _next_reg_T_37 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1436 = 5'h1b == rd ? _next_reg_T_37 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1437 = 5'h1c == rd ? _next_reg_T_37 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1438 = 5'h1d == rd ? _next_reg_T_37 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1439 = 5'h1e == rd ? _next_reg_T_37 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1440 = 5'h1f == rd ? _next_reg_T_37 : _GEN_1408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [6:0] _GEN_1442 = _T_119 ? inst[31:25] : _GEN_1371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1445 = _T_119 ? inst[14:12] : _GEN_1374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1447 = _T_119 ? inst[6:0] : _GEN_1376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1448 = _T_119 ? _GEN_1409 : _GEN_1377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1449 = _T_119 ? _GEN_1410 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1450 = _T_119 ? _GEN_1411 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1451 = _T_119 ? _GEN_1412 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1452 = _T_119 ? _GEN_1413 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1453 = _T_119 ? _GEN_1414 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1454 = _T_119 ? _GEN_1415 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1455 = _T_119 ? _GEN_1416 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1456 = _T_119 ? _GEN_1417 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1457 = _T_119 ? _GEN_1418 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1458 = _T_119 ? _GEN_1419 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1459 = _T_119 ? _GEN_1420 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1460 = _T_119 ? _GEN_1421 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1461 = _T_119 ? _GEN_1422 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1462 = _T_119 ? _GEN_1423 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1463 = _T_119 ? _GEN_1424 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1464 = _T_119 ? _GEN_1425 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1465 = _T_119 ? _GEN_1426 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1466 = _T_119 ? _GEN_1427 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1467 = _T_119 ? _GEN_1428 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1468 = _T_119 ? _GEN_1429 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1469 = _T_119 ? _GEN_1430 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1470 = _T_119 ? _GEN_1431 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1471 = _T_119 ? _GEN_1432 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1472 = _T_119 ? _GEN_1433 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1473 = _T_119 ? _GEN_1434 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1474 = _T_119 ? _GEN_1435 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1475 = _T_119 ? _GEN_1436 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1476 = _T_119 ? _GEN_1437 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1477 = _T_119 ? _GEN_1438 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1478 = _T_119 ? _GEN_1439 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1479 = _T_119 ? _GEN_1440 : _GEN_1408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [6:0] _funct7_T_9 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_18 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_131 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_17 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_38 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:62]
  wire [31:0] _now_reg_rs2_8 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [4:0] _next_reg_T_39 = _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:84]
  wire [31:0] _next_reg_T_40 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:69]
  wire [31:0] _next_reg_T_41 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:92]
  wire [31:0] _next_reg_rd_19 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:92]
  wire [31:0] _GEN_1480 = 5'h0 == rd ? _next_reg_T_41 : _GEN_1448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1481 = 5'h1 == rd ? _next_reg_T_41 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1482 = 5'h2 == rd ? _next_reg_T_41 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1483 = 5'h3 == rd ? _next_reg_T_41 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1484 = 5'h4 == rd ? _next_reg_T_41 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1485 = 5'h5 == rd ? _next_reg_T_41 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1486 = 5'h6 == rd ? _next_reg_T_41 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1487 = 5'h7 == rd ? _next_reg_T_41 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1488 = 5'h8 == rd ? _next_reg_T_41 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1489 = 5'h9 == rd ? _next_reg_T_41 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1490 = 5'ha == rd ? _next_reg_T_41 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1491 = 5'hb == rd ? _next_reg_T_41 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1492 = 5'hc == rd ? _next_reg_T_41 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1493 = 5'hd == rd ? _next_reg_T_41 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1494 = 5'he == rd ? _next_reg_T_41 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1495 = 5'hf == rd ? _next_reg_T_41 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1496 = 5'h10 == rd ? _next_reg_T_41 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1497 = 5'h11 == rd ? _next_reg_T_41 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1498 = 5'h12 == rd ? _next_reg_T_41 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1499 = 5'h13 == rd ? _next_reg_T_41 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1500 = 5'h14 == rd ? _next_reg_T_41 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1501 = 5'h15 == rd ? _next_reg_T_41 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1502 = 5'h16 == rd ? _next_reg_T_41 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1503 = 5'h17 == rd ? _next_reg_T_41 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1504 = 5'h18 == rd ? _next_reg_T_41 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1505 = 5'h19 == rd ? _next_reg_T_41 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1506 = 5'h1a == rd ? _next_reg_T_41 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1507 = 5'h1b == rd ? _next_reg_T_41 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1508 = 5'h1c == rd ? _next_reg_T_41 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1509 = 5'h1d == rd ? _next_reg_T_41 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1510 = 5'h1e == rd ? _next_reg_T_41 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1511 = 5'h1f == rd ? _next_reg_T_41 : _GEN_1479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [6:0] _GEN_1513 = _T_126 ? inst[31:25] : _GEN_1442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1516 = _T_126 ? inst[14:12] : _GEN_1445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1518 = _T_126 ? inst[6:0] : _GEN_1447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1519 = _T_126 ? _GEN_1480 : _GEN_1448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1520 = _T_126 ? _GEN_1481 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1521 = _T_126 ? _GEN_1482 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1522 = _T_126 ? _GEN_1483 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1523 = _T_126 ? _GEN_1484 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1524 = _T_126 ? _GEN_1485 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1525 = _T_126 ? _GEN_1486 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1526 = _T_126 ? _GEN_1487 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1527 = _T_126 ? _GEN_1488 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1528 = _T_126 ? _GEN_1489 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1529 = _T_126 ? _GEN_1490 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1530 = _T_126 ? _GEN_1491 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1531 = _T_126 ? _GEN_1492 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1532 = _T_126 ? _GEN_1493 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1533 = _T_126 ? _GEN_1494 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1534 = _T_126 ? _GEN_1495 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1535 = _T_126 ? _GEN_1496 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1536 = _T_126 ? _GEN_1497 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1537 = _T_126 ? _GEN_1498 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1538 = _T_126 ? _GEN_1499 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1539 = _T_126 ? _GEN_1500 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1540 = _T_126 ? _GEN_1501 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1541 = _T_126 ? _GEN_1502 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1542 = _T_126 ? _GEN_1503 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1543 = _T_126 ? _GEN_1504 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1544 = _T_126 ? _GEN_1505 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1545 = _T_126 ? _GEN_1506 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1546 = _T_126 ? _GEN_1507 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1547 = _T_126 ? _GEN_1508 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1548 = _T_126 ? _GEN_1509 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1549 = _T_126 ? _GEN_1510 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1550 = _T_126 ? _GEN_1511 : _GEN_1479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [6:0] _T_138 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 191:37]
  wire [31:0] _next_pc_T_1 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 191:37]
  wire [32:0] _next_reg_T_42 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [31:0] _next_reg_T_43 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [31:0] _next_reg_rd_20 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [31:0] _GEN_1551 = 5'h0 == rd ? _next_reg_T_43 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1552 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1553 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1554 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1555 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1556 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1557 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1558 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1559 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1560 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1561 = 5'ha == rd ? _next_reg_T_43 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1562 = 5'hb == rd ? _next_reg_T_43 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1563 = 5'hc == rd ? _next_reg_T_43 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1564 = 5'hd == rd ? _next_reg_T_43 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1565 = 5'he == rd ? _next_reg_T_43 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1566 = 5'hf == rd ? _next_reg_T_43 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1567 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1568 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1569 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1570 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1571 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1572 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1573 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1574 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1575 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1576 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1577 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1578 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1579 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1580 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1581 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1582 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [32:0] _next_csr_mtval_T = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 194:34]
  wire [31:0] _next_csr_mtval_T_1 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 194:34]
  wire  _GEN_1583 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _GEN_1584 = _T_346 ? _T_334 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 191:27]
  wire [31:0] _GEN_1585 = _T_346 ? _GEN_1551 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1586 = _T_346 ? _GEN_1552 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1587 = _T_346 ? _GEN_1553 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1588 = _T_346 ? _GEN_1554 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1589 = _T_346 ? _GEN_1555 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1590 = _T_346 ? _GEN_1556 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1591 = _T_346 ? _GEN_1557 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1592 = _T_346 ? _GEN_1558 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1593 = _T_346 ? _GEN_1559 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1594 = _T_346 ? _GEN_1560 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1595 = _T_346 ? _GEN_1561 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1596 = _T_346 ? _GEN_1562 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1597 = _T_346 ? _GEN_1563 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1598 = _T_346 ? _GEN_1564 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1599 = _T_346 ? _GEN_1565 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1600 = _T_346 ? _GEN_1566 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1601 = _T_346 ? _GEN_1567 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1602 = _T_346 ? _GEN_1568 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1603 = _T_346 ? _GEN_1569 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1604 = _T_346 ? _GEN_1570 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1605 = _T_346 ? _GEN_1571 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1606 = _T_346 ? _GEN_1572 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1607 = _T_346 ? _GEN_1573 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1608 = _T_346 ? _GEN_1574 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1609 = _T_346 ? _GEN_1575 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1610 = _T_346 ? _GEN_1576 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1611 = _T_346 ? _GEN_1577 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1612 = _T_346 ? _GEN_1578 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1613 = _T_346 ? _GEN_1579 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1614 = _T_346 ? _GEN_1580 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1615 = _T_346 ? _GEN_1581 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1616 = _T_346 ? _GEN_1582 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] now_csr_mtval = io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_1617 = _T_346 ? io_now_csr_mtval : _T_334; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 194:24]
  wire  _GEN_1619 = _T_346 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36 145:33]
  wire [6:0] _GEN_1626 = _T_133 ? inst[6:0] : _GEN_1518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1628 = _T_133 & _T_346; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 113:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1629 = _T_133 ? _GEN_1584 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1630 = _T_133 ? _GEN_1585 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1631 = _T_133 ? _GEN_1586 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1632 = _T_133 ? _GEN_1587 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1633 = _T_133 ? _GEN_1588 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1634 = _T_133 ? _GEN_1589 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1635 = _T_133 ? _GEN_1590 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1636 = _T_133 ? _GEN_1591 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1637 = _T_133 ? _GEN_1592 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1638 = _T_133 ? _GEN_1593 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1639 = _T_133 ? _GEN_1594 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1640 = _T_133 ? _GEN_1595 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1641 = _T_133 ? _GEN_1596 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1642 = _T_133 ? _GEN_1597 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1643 = _T_133 ? _GEN_1598 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1644 = _T_133 ? _GEN_1599 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1645 = _T_133 ? _GEN_1600 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1646 = _T_133 ? _GEN_1601 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1647 = _T_133 ? _GEN_1602 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1648 = _T_133 ? _GEN_1603 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1649 = _T_133 ? _GEN_1604 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1650 = _T_133 ? _GEN_1605 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1651 = _T_133 ? _GEN_1606 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1652 = _T_133 ? _GEN_1607 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1653 = _T_133 ? _GEN_1608 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1654 = _T_133 ? _GEN_1609 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1655 = _T_133 ? _GEN_1610 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1656 = _T_133 ? _GEN_1611 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1657 = _T_133 ? _GEN_1612 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1658 = _T_133 ? _GEN_1613 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1659 = _T_133 ? _GEN_1614 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1660 = _T_133 ? _GEN_1615 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1661 = _T_133 ? _GEN_1616 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1662 = _T_133 ? _GEN_1617 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire  _GEN_1664 = _T_133 & _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [2:0] _funct3_T_19 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_161 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_19 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_pc_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:48]
  wire [31:0] _next_pc_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:48]
  wire [30:0] _next_pc_T_4 = _T_433[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:54]
  wire [31:0] _next_pc_T_5 = {_T_433[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:33]
  wire [32:0] _next_reg_T_44 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:37]
  wire [31:0] _next_reg_T_45 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:37]
  wire [31:0] _next_reg_rd_21 = _next_reg_T_43; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:37]
  wire [31:0] _GEN_1665 = 5'h0 == rd ? _next_reg_T_43 : _GEN_1630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1666 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1667 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1668 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1669 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1670 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1671 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1672 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1673 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1674 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1675 = 5'ha == rd ? _next_reg_T_43 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1676 = 5'hb == rd ? _next_reg_T_43 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1677 = 5'hc == rd ? _next_reg_T_43 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1678 = 5'hd == rd ? _next_reg_T_43 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1679 = 5'he == rd ? _next_reg_T_43 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1680 = 5'hf == rd ? _next_reg_T_43 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1681 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1682 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1683 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1684 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1685 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1686 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1687 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1688 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1689 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1690 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1691 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1692 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1693 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1694 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1695 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1696 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _now_reg_rs1_20 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_csr_mtval_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:45]
  wire [31:0] _next_csr_mtval_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:45]
  wire [30:0] _next_csr_mtval_T_4 = _T_433[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:51]
  wire [31:0] _next_csr_mtval_T_5 = {_T_433[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:30]
  wire  _GEN_1697 = _T_180 | _GEN_1628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 202:27]
  wire [31:0] _GEN_1698 = _T_180 ? _T_168 : _GEN_1629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 203:27]
  wire [31:0] _GEN_1699 = _T_180 ? _GEN_1665 : _GEN_1630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1700 = _T_180 ? _GEN_1666 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1701 = _T_180 ? _GEN_1667 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1702 = _T_180 ? _GEN_1668 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1703 = _T_180 ? _GEN_1669 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1704 = _T_180 ? _GEN_1670 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1705 = _T_180 ? _GEN_1671 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1706 = _T_180 ? _GEN_1672 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1707 = _T_180 ? _GEN_1673 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1708 = _T_180 ? _GEN_1674 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1709 = _T_180 ? _GEN_1675 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1710 = _T_180 ? _GEN_1676 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1711 = _T_180 ? _GEN_1677 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1712 = _T_180 ? _GEN_1678 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1713 = _T_180 ? _GEN_1679 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1714 = _T_180 ? _GEN_1680 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1715 = _T_180 ? _GEN_1681 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1716 = _T_180 ? _GEN_1682 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1717 = _T_180 ? _GEN_1683 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1718 = _T_180 ? _GEN_1684 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1719 = _T_180 ? _GEN_1685 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1720 = _T_180 ? _GEN_1686 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1721 = _T_180 ? _GEN_1687 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1722 = _T_180 ? _GEN_1688 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1723 = _T_180 ? _GEN_1689 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1724 = _T_180 ? _GEN_1690 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1725 = _T_180 ? _GEN_1691 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1726 = _T_180 ? _GEN_1692 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1727 = _T_180 ? _GEN_1693 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1728 = _T_180 ? _GEN_1694 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1729 = _T_180 ? _GEN_1695 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1730 = _T_180 ? _GEN_1696 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1731 = _T_180 ? _GEN_1662 : _T_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 206:24]
  wire  _GEN_1733 = _T_180 ? _GEN_1663 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_1737 = _T_157 ? inst[14:12] : _GEN_1516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1739 = _T_157 ? inst[6:0] : _GEN_1626; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1741 = _T_157 ? _GEN_1697 : _GEN_1628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1742 = _T_157 ? _GEN_1698 : _GEN_1629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1743 = _T_157 ? _GEN_1699 : _GEN_1630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1744 = _T_157 ? _GEN_1700 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1745 = _T_157 ? _GEN_1701 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1746 = _T_157 ? _GEN_1702 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1747 = _T_157 ? _GEN_1703 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1748 = _T_157 ? _GEN_1704 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1749 = _T_157 ? _GEN_1705 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1750 = _T_157 ? _GEN_1706 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1751 = _T_157 ? _GEN_1707 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1752 = _T_157 ? _GEN_1708 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1753 = _T_157 ? _GEN_1709 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1754 = _T_157 ? _GEN_1710 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1755 = _T_157 ? _GEN_1711 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1756 = _T_157 ? _GEN_1712 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1757 = _T_157 ? _GEN_1713 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1758 = _T_157 ? _GEN_1714 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1759 = _T_157 ? _GEN_1715 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1760 = _T_157 ? _GEN_1716 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1761 = _T_157 ? _GEN_1717 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1762 = _T_157 ? _GEN_1718 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1763 = _T_157 ? _GEN_1719 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1764 = _T_157 ? _GEN_1720 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1765 = _T_157 ? _GEN_1721 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1766 = _T_157 ? _GEN_1722 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1767 = _T_157 ? _GEN_1723 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1768 = _T_157 ? _GEN_1724 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1769 = _T_157 ? _GEN_1725 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1770 = _T_157 ? _GEN_1726 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1771 = _T_157 ? _GEN_1727 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1772 = _T_157 ? _GEN_1728 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1773 = _T_157 ? _GEN_1729 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1774 = _T_157 ? _GEN_1730 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1775 = _T_157 ? _GEN_1731 : _GEN_1662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1777 = _T_157 ? _GEN_1732 : _GEN_1663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [2:0] _funct3_T_20 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_189 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_6 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 217:39]
  wire [31:0] _next_pc_T_7 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 217:39]
  wire [32:0] _next_csr_mtval_T_6 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 219:36]
  wire [31:0] _next_csr_mtval_T_7 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 219:36]
  wire  _GEN_1778 = _T_346 | _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 216:29]
  wire [31:0] _GEN_1779 = _T_346 ? _T_334 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 217:29]
  wire [31:0] _GEN_1780 = _T_346 ? _GEN_1775 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 219:26]
  wire  _GEN_1782 = _T_346 ? _GEN_1776 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1783 = _GEN_31 == _GEN_840 ? _GEN_1778 : _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [31:0] _GEN_1784 = _GEN_31 == _GEN_840 ? _GEN_1779 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [31:0] _GEN_1785 = _GEN_31 == _GEN_840 ? _GEN_1780 : _GEN_1775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1787 = _GEN_31 == _GEN_840 ? _GEN_1781 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [2:0] _GEN_1793 = _T_182 ? inst[14:12] : _GEN_1737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1796 = _T_182 ? inst[6:0] : _GEN_1739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1798 = _T_182 ? _GEN_1783 : _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [31:0] _GEN_1799 = _T_182 ? _GEN_1784 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [31:0] _GEN_1800 = _T_182 ? _GEN_1785 : _GEN_1775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1802 = _T_182 ? _GEN_1786 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [2:0] _funct3_T_21 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_216 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_8 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 229:39]
  wire [31:0] _next_pc_T_9 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 229:39]
  wire [32:0] _next_csr_mtval_T_8 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 231:36]
  wire [31:0] _next_csr_mtval_T_9 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 231:36]
  wire  _GEN_1803 = _T_346 | _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 228:29]
  wire [31:0] _GEN_1804 = _T_346 ? _T_334 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 229:29]
  wire [31:0] _GEN_1805 = _T_346 ? _GEN_1800 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 231:26]
  wire  _GEN_1807 = _T_346 ? _GEN_1801 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1808 = _GEN_31 != _GEN_840 ? _GEN_1803 : _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [31:0] _GEN_1809 = _GEN_31 != _GEN_840 ? _GEN_1804 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [31:0] _GEN_1810 = _GEN_31 != _GEN_840 ? _GEN_1805 : _GEN_1800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1812 = _GEN_31 != _GEN_840 ? _GEN_1806 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [2:0] _GEN_1818 = _T_209 ? inst[14:12] : _GEN_1793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1821 = _T_209 ? inst[6:0] : _GEN_1796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1823 = _T_209 ? _GEN_1808 : _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [31:0] _GEN_1824 = _T_209 ? _GEN_1809 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [31:0] _GEN_1825 = _T_209 ? _GEN_1810 : _GEN_1800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1827 = _T_209 ? _GEN_1811 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [2:0] _funct3_T_22 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_243 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_10 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 242:39]
  wire [31:0] _next_pc_T_11 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 242:39]
  wire [32:0] _next_csr_mtval_T_10 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 244:36]
  wire [31:0] _next_csr_mtval_T_11 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 244:36]
  wire  _GEN_1828 = _T_346 | _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 241:29]
  wire [31:0] _GEN_1829 = _T_346 ? _T_334 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 242:29]
  wire [31:0] _GEN_1830 = _T_346 ? _GEN_1825 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 244:26]
  wire  _GEN_1832 = _T_346 ? _GEN_1826 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1833 = $signed(_T_300) < $signed(_T_301) ? _GEN_1828 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [31:0] _GEN_1834 = $signed(_T_300) < $signed(_T_301) ? _GEN_1829 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [31:0] _GEN_1835 = $signed(_T_300) < $signed(_T_301) ? _GEN_1830 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1837 = $signed(_T_300) < $signed(_T_301) ? _GEN_1831 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [2:0] _GEN_1843 = _T_236 ? inst[14:12] : _GEN_1818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1846 = _T_236 ? inst[6:0] : _GEN_1821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1848 = _T_236 ? _GEN_1833 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [31:0] _GEN_1849 = _T_236 ? _GEN_1834 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [31:0] _GEN_1850 = _T_236 ? _GEN_1835 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1852 = _T_236 ? _GEN_1836 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [2:0] _funct3_T_23 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_272 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_12 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 254:39]
  wire [31:0] _next_pc_T_13 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 254:39]
  wire [32:0] _next_csr_mtval_T_12 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 256:36]
  wire [31:0] _next_csr_mtval_T_13 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 256:36]
  wire  _GEN_1853 = _T_346 | _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 253:29]
  wire [31:0] _GEN_1854 = _T_346 ? _T_334 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 254:29]
  wire [31:0] _GEN_1855 = _T_346 ? _GEN_1850 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 256:26]
  wire  _GEN_1857 = _T_346 ? _GEN_1851 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1858 = _GEN_31 < _GEN_840 ? _GEN_1853 : _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [31:0] _GEN_1859 = _GEN_31 < _GEN_840 ? _GEN_1854 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [31:0] _GEN_1860 = _GEN_31 < _GEN_840 ? _GEN_1855 : _GEN_1850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1862 = _GEN_31 < _GEN_840 ? _GEN_1856 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [2:0] _GEN_1868 = _T_265 ? inst[14:12] : _GEN_1843; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1871 = _T_265 ? inst[6:0] : _GEN_1846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1873 = _T_265 ? _GEN_1858 : _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [31:0] _GEN_1874 = _T_265 ? _GEN_1859 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [31:0] _GEN_1875 = _T_265 ? _GEN_1860 : _GEN_1850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1877 = _T_265 ? _GEN_1861 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [2:0] _funct3_T_24 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_299 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_14 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 267:39]
  wire [31:0] _next_pc_T_15 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 267:39]
  wire [32:0] _next_csr_mtval_T_14 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 269:36]
  wire [31:0] _next_csr_mtval_T_15 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 269:36]
  wire  _GEN_1878 = _T_346 | _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 266:29]
  wire [31:0] _GEN_1879 = _T_346 ? _T_334 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 267:29]
  wire [31:0] _GEN_1880 = _T_346 ? _GEN_1875 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 269:26]
  wire  _GEN_1882 = _T_346 ? _GEN_1876 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1883 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1878 : _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [31:0] _GEN_1884 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1879 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [31:0] _GEN_1885 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1880 : _GEN_1875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1887 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1881 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [2:0] _GEN_1893 = _T_292 ? inst[14:12] : _GEN_1868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1896 = _T_292 ? inst[6:0] : _GEN_1871; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1898 = _T_292 ? _GEN_1883 : _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [31:0] _GEN_1899 = _T_292 ? _GEN_1884 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [31:0] _GEN_1900 = _T_292 ? _GEN_1885 : _GEN_1875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1902 = _T_292 ? _GEN_1886 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [2:0] _funct3_T_25 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_328 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_16 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 279:39]
  wire [31:0] _next_pc_T_17 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 279:39]
  wire [32:0] _next_csr_mtval_T_16 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 281:36]
  wire [31:0] _next_csr_mtval_T_17 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 281:36]
  wire  _GEN_1903 = _T_346 | _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 278:29]
  wire [31:0] _GEN_1904 = _T_346 ? _T_334 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 279:29]
  wire [31:0] _GEN_1905 = _T_346 ? _GEN_1900 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 281:26]
  wire  _GEN_1907 = _T_346 ? _GEN_1901 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1908 = _GEN_31 >= _GEN_840 ? _GEN_1903 : _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [31:0] _GEN_1909 = _GEN_31 >= _GEN_840 ? _GEN_1904 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [31:0] _GEN_1910 = _GEN_31 >= _GEN_840 ? _GEN_1905 : _GEN_1900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1912 = _GEN_31 >= _GEN_840 ? _GEN_1906 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [2:0] _GEN_1918 = _T_321 ? inst[14:12] : _GEN_1893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1921 = _T_321 ? inst[6:0] : _GEN_1896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1923 = _T_321 ? _GEN_1908 : _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [31:0] _GEN_1924 = _T_321 ? _GEN_1909 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [31:0] _GEN_1925 = _T_321 ? _GEN_1910 : _GEN_1900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  _GEN_1927 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [2:0] _funct3_T_26 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_352 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_28 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_46 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:54]
  wire [31:0] _next_reg_T_47 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:54]
  wire [1:0] _next_reg_rOff_T = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_1 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_2 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_3 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_4 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_5 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_6 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 164:10 21:22]
  wire [31:0] _next_reg_T_48 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6207 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_49 = _GEN_6207 & 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [7:0] _next_reg_T_50 = _next_reg_T_49[7:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:65]
  wire  next_reg_signBit = _next_reg_T_49[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _next_reg_T_51 = next_reg_signBit; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [23:0] _next_reg_T_52 = next_reg_signBit ? 24'hffffff : 24'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _next_reg_T_53 = {_next_reg_T_52,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _next_reg_rd_22 = {_next_reg_T_52,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_1928 = 5'h0 == rd ? _next_reg_T_53 : _GEN_1743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1929 = 5'h1 == rd ? _next_reg_T_53 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1930 = 5'h2 == rd ? _next_reg_T_53 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1931 = 5'h3 == rd ? _next_reg_T_53 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1932 = 5'h4 == rd ? _next_reg_T_53 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1933 = 5'h5 == rd ? _next_reg_T_53 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1934 = 5'h6 == rd ? _next_reg_T_53 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1935 = 5'h7 == rd ? _next_reg_T_53 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1936 = 5'h8 == rd ? _next_reg_T_53 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1937 = 5'h9 == rd ? _next_reg_T_53 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1938 = 5'ha == rd ? _next_reg_T_53 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1939 = 5'hb == rd ? _next_reg_T_53 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1940 = 5'hc == rd ? _next_reg_T_53 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1941 = 5'hd == rd ? _next_reg_T_53 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1942 = 5'he == rd ? _next_reg_T_53 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1943 = 5'hf == rd ? _next_reg_T_53 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1944 = 5'h10 == rd ? _next_reg_T_53 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1945 = 5'h11 == rd ? _next_reg_T_53 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1946 = 5'h12 == rd ? _next_reg_T_53 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1947 = 5'h13 == rd ? _next_reg_T_53 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1948 = 5'h14 == rd ? _next_reg_T_53 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1949 = 5'h15 == rd ? _next_reg_T_53 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1950 = 5'h16 == rd ? _next_reg_T_53 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1951 = 5'h17 == rd ? _next_reg_T_53 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1952 = 5'h18 == rd ? _next_reg_T_53 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1953 = 5'h19 == rd ? _next_reg_T_53 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1954 = 5'h1a == rd ? _next_reg_T_53 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1955 = 5'h1b == rd ? _next_reg_T_53 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1956 = 5'h1c == rd ? _next_reg_T_53 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1957 = 5'h1d == rd ? _next_reg_T_53 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1958 = 5'h1e == rd ? _next_reg_T_53 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1959 = 5'h1f == rd ? _next_reg_T_53 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _now_reg_rs1_29 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 294:39]
  wire [31:0] _mem_read_addr_T_1 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 294:39]
  wire  _mem_WIRE_read_valid = 1'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire  _GEN_1960 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _GEN_1961 = _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:54]
  wire [5:0] _mem_WIRE_read_memWidth = 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [5:0] _GEN_1962 = 6'h8; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _GEN_1963 = 5'h0 == rd ? _next_reg_T_53 : _GEN_1743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1964 = 5'h1 == rd ? _next_reg_T_53 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1965 = 5'h2 == rd ? _next_reg_T_53 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1966 = 5'h3 == rd ? _next_reg_T_53 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1967 = 5'h4 == rd ? _next_reg_T_53 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1968 = 5'h5 == rd ? _next_reg_T_53 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1969 = 5'h6 == rd ? _next_reg_T_53 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1970 = 5'h7 == rd ? _next_reg_T_53 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1971 = 5'h8 == rd ? _next_reg_T_53 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1972 = 5'h9 == rd ? _next_reg_T_53 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1973 = 5'ha == rd ? _next_reg_T_53 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1974 = 5'hb == rd ? _next_reg_T_53 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1975 = 5'hc == rd ? _next_reg_T_53 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1976 = 5'hd == rd ? _next_reg_T_53 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1977 = 5'he == rd ? _next_reg_T_53 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1978 = 5'hf == rd ? _next_reg_T_53 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1979 = 5'h10 == rd ? _next_reg_T_53 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1980 = 5'h11 == rd ? _next_reg_T_53 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1981 = 5'h12 == rd ? _next_reg_T_53 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1982 = 5'h13 == rd ? _next_reg_T_53 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1983 = 5'h14 == rd ? _next_reg_T_53 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1984 = 5'h15 == rd ? _next_reg_T_53 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1985 = 5'h16 == rd ? _next_reg_T_53 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1986 = 5'h17 == rd ? _next_reg_T_53 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1987 = 5'h18 == rd ? _next_reg_T_53 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1988 = 5'h19 == rd ? _next_reg_T_53 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1989 = 5'h1a == rd ? _next_reg_T_53 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1990 = 5'h1b == rd ? _next_reg_T_53 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1991 = 5'h1c == rd ? _next_reg_T_53 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1992 = 5'h1d == rd ? _next_reg_T_53 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1993 = 5'h1e == rd ? _next_reg_T_53 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1994 = 5'h1f == rd ? _next_reg_T_53 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire  _GEN_1996 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [2:0] _GEN_2000 = _T_348 ? inst[14:12] : _GEN_1918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2002 = _T_348 ? inst[6:0] : _GEN_1921; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2004 = 32'h3 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _mem_WIRE_read_addr = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [31:0] _GEN_2005 = _T_348 ? _T_433 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [5:0] _GEN_2006 = _T_348 ? 6'h8 : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _GEN_2007 = _T_348 ? _GEN_1928 : _GEN_1743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2008 = _T_348 ? _GEN_1929 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2009 = _T_348 ? _GEN_1930 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2010 = _T_348 ? _GEN_1931 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2011 = _T_348 ? _GEN_1932 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2012 = _T_348 ? _GEN_1933 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2013 = _T_348 ? _GEN_1934 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2014 = _T_348 ? _GEN_1935 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2015 = _T_348 ? _GEN_1936 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2016 = _T_348 ? _GEN_1937 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2017 = _T_348 ? _GEN_1938 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2018 = _T_348 ? _GEN_1939 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2019 = _T_348 ? _GEN_1940 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2020 = _T_348 ? _GEN_1941 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2021 = _T_348 ? _GEN_1942 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2022 = _T_348 ? _GEN_1943 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2023 = _T_348 ? _GEN_1944 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2024 = _T_348 ? _GEN_1945 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2025 = _T_348 ? _GEN_1946 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2026 = _T_348 ? _GEN_1947 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2027 = _T_348 ? _GEN_1948 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2028 = _T_348 ? _GEN_1949 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2029 = _T_348 ? _GEN_1950 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2030 = _T_348 ? _GEN_1951 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2031 = _T_348 ? _GEN_1952 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2032 = _T_348 ? _GEN_1953 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2033 = _T_348 ? _GEN_1954 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2034 = _T_348 ? _GEN_1955 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2035 = _T_348 ? _GEN_1956 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2036 = _T_348 ? _GEN_1957 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2037 = _T_348 ? _GEN_1958 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2038 = _T_348 ? _GEN_1959 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire  _GEN_2040 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [2:0] _funct3_T_27 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_372 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_31 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_54 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:54]
  wire [31:0] _next_reg_T_55 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:54]
  wire [1:0] _next_reg_rOff_T_1 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_1 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_7 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_8 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_9 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_10 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_11 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_12 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_13 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_1 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_56 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6208 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_57 = _GEN_6207 & 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [15:0] _next_reg_T_58 = _next_reg_T_57[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:66]
  wire  next_reg_signBit_1 = _next_reg_T_57[15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _next_reg_T_59 = next_reg_signBit_1; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [15:0] _next_reg_T_60 = next_reg_signBit_1 ? 16'hffff : 16'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _next_reg_T_61 = {_next_reg_T_60,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _next_reg_rd_23 = {_next_reg_T_60,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_2041 = 5'h0 == rd ? _next_reg_T_61 : _GEN_2007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2042 = 5'h1 == rd ? _next_reg_T_61 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2043 = 5'h2 == rd ? _next_reg_T_61 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2044 = 5'h3 == rd ? _next_reg_T_61 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2045 = 5'h4 == rd ? _next_reg_T_61 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2046 = 5'h5 == rd ? _next_reg_T_61 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2047 = 5'h6 == rd ? _next_reg_T_61 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2048 = 5'h7 == rd ? _next_reg_T_61 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2049 = 5'h8 == rd ? _next_reg_T_61 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2050 = 5'h9 == rd ? _next_reg_T_61 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2051 = 5'ha == rd ? _next_reg_T_61 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2052 = 5'hb == rd ? _next_reg_T_61 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2053 = 5'hc == rd ? _next_reg_T_61 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2054 = 5'hd == rd ? _next_reg_T_61 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2055 = 5'he == rd ? _next_reg_T_61 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2056 = 5'hf == rd ? _next_reg_T_61 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2057 = 5'h10 == rd ? _next_reg_T_61 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2058 = 5'h11 == rd ? _next_reg_T_61 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2059 = 5'h12 == rd ? _next_reg_T_61 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2060 = 5'h13 == rd ? _next_reg_T_61 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2061 = 5'h14 == rd ? _next_reg_T_61 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2062 = 5'h15 == rd ? _next_reg_T_61 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2063 = 5'h16 == rd ? _next_reg_T_61 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2064 = 5'h17 == rd ? _next_reg_T_61 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2065 = 5'h18 == rd ? _next_reg_T_61 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2066 = 5'h19 == rd ? _next_reg_T_61 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2067 = 5'h1a == rd ? _next_reg_T_61 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2068 = 5'h1b == rd ? _next_reg_T_61 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2069 = 5'h1c == rd ? _next_reg_T_61 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2070 = 5'h1d == rd ? _next_reg_T_61 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2071 = 5'h1e == rd ? _next_reg_T_61 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2072 = 5'h1f == rd ? _next_reg_T_61 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _now_reg_rs1_32 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 303:39]
  wire [31:0] _mem_read_addr_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 303:39]
  wire  _GEN_2073 = _T_435 | _T_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2074 = _T_435 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 303:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2075 = _T_435 ? 6'h10 : _GEN_2006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2076 = _T_435 ? _GEN_2041 : _GEN_2007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2077 = _T_435 ? _GEN_2042 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2078 = _T_435 ? _GEN_2043 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2079 = _T_435 ? _GEN_2044 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2080 = _T_435 ? _GEN_2045 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2081 = _T_435 ? _GEN_2046 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2082 = _T_435 ? _GEN_2047 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2083 = _T_435 ? _GEN_2048 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2084 = _T_435 ? _GEN_2049 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2085 = _T_435 ? _GEN_2050 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2086 = _T_435 ? _GEN_2051 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2087 = _T_435 ? _GEN_2052 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2088 = _T_435 ? _GEN_2053 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2089 = _T_435 ? _GEN_2054 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2090 = _T_435 ? _GEN_2055 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2091 = _T_435 ? _GEN_2056 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2092 = _T_435 ? _GEN_2057 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2093 = _T_435 ? _GEN_2058 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2094 = _T_435 ? _GEN_2059 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2095 = _T_435 ? _GEN_2060 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2096 = _T_435 ? _GEN_2061 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2097 = _T_435 ? _GEN_2062 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2098 = _T_435 ? _GEN_2063 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2099 = _T_435 ? _GEN_2064 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2100 = _T_435 ? _GEN_2065 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2101 = _T_435 ? _GEN_2066 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2102 = _T_435 ? _GEN_2067 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2103 = _T_435 ? _GEN_2068 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2104 = _T_435 ? _GEN_2069 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2105 = _T_435 ? _GEN_2070 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2106 = _T_435 ? _GEN_2071 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2107 = _T_435 ? _GEN_2072 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2109 = _T_435 ? _GEN_1926 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2113 = _T_368 ? inst[14:12] : _GEN_2000; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2115 = _T_368 ? inst[6:0] : _GEN_2002; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2117 = _T_368 ? _GEN_2073 : _T_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2118 = _T_368 ? _GEN_2074 : _GEN_2005; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [5:0] _GEN_2119 = _T_368 ? _GEN_2075 : _GEN_2006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2120 = _T_368 ? _GEN_2076 : _GEN_2007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2121 = _T_368 ? _GEN_2077 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2122 = _T_368 ? _GEN_2078 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2123 = _T_368 ? _GEN_2079 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2124 = _T_368 ? _GEN_2080 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2125 = _T_368 ? _GEN_2081 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2126 = _T_368 ? _GEN_2082 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2127 = _T_368 ? _GEN_2083 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2128 = _T_368 ? _GEN_2084 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2129 = _T_368 ? _GEN_2085 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2130 = _T_368 ? _GEN_2086 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2131 = _T_368 ? _GEN_2087 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2132 = _T_368 ? _GEN_2088 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2133 = _T_368 ? _GEN_2089 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2134 = _T_368 ? _GEN_2090 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2135 = _T_368 ? _GEN_2091 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2136 = _T_368 ? _GEN_2092 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2137 = _T_368 ? _GEN_2093 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2138 = _T_368 ? _GEN_2094 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2139 = _T_368 ? _GEN_2095 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2140 = _T_368 ? _GEN_2096 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2141 = _T_368 ? _GEN_2097 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2142 = _T_368 ? _GEN_2098 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2143 = _T_368 ? _GEN_2099 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2144 = _T_368 ? _GEN_2100 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2145 = _T_368 ? _GEN_2101 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2146 = _T_368 ? _GEN_2102 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2147 = _T_368 ? _GEN_2103 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2148 = _T_368 ? _GEN_2104 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2149 = _T_368 ? _GEN_2105 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2150 = _T_368 ? _GEN_2106 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2151 = _T_368 ? _GEN_2107 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2153 = _T_368 ? _GEN_2109 : _GEN_1926; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [2:0] _funct3_T_28 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_392 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_34 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_62 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:54]
  wire [31:0] _next_reg_T_63 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:54]
  wire [1:0] _next_reg_rOff_T_2 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_2 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_14 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_15 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_16 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_17 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_18 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_19 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_20 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_2 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_64 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6209 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_65 = _GEN_6207 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [31:0] _next_reg_T_66 = _next_reg_T_65[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:66]
  wire  next_reg_signBit_2 = _next_reg_T_65[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_67 = _next_reg_T_65[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:66]
  wire [31:0] _next_reg_rd_24 = _next_reg_T_65[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:66]
  wire [31:0] _GEN_2154 = 5'h0 == rd ? _next_reg_T_65[31:0] : _GEN_2120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2155 = 5'h1 == rd ? _next_reg_T_65[31:0] : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2156 = 5'h2 == rd ? _next_reg_T_65[31:0] : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2157 = 5'h3 == rd ? _next_reg_T_65[31:0] : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2158 = 5'h4 == rd ? _next_reg_T_65[31:0] : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2159 = 5'h5 == rd ? _next_reg_T_65[31:0] : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2160 = 5'h6 == rd ? _next_reg_T_65[31:0] : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2161 = 5'h7 == rd ? _next_reg_T_65[31:0] : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2162 = 5'h8 == rd ? _next_reg_T_65[31:0] : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2163 = 5'h9 == rd ? _next_reg_T_65[31:0] : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2164 = 5'ha == rd ? _next_reg_T_65[31:0] : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2165 = 5'hb == rd ? _next_reg_T_65[31:0] : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2166 = 5'hc == rd ? _next_reg_T_65[31:0] : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2167 = 5'hd == rd ? _next_reg_T_65[31:0] : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2168 = 5'he == rd ? _next_reg_T_65[31:0] : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2169 = 5'hf == rd ? _next_reg_T_65[31:0] : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2170 = 5'h10 == rd ? _next_reg_T_65[31:0] : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2171 = 5'h11 == rd ? _next_reg_T_65[31:0] : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2172 = 5'h12 == rd ? _next_reg_T_65[31:0] : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2173 = 5'h13 == rd ? _next_reg_T_65[31:0] : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2174 = 5'h14 == rd ? _next_reg_T_65[31:0] : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2175 = 5'h15 == rd ? _next_reg_T_65[31:0] : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2176 = 5'h16 == rd ? _next_reg_T_65[31:0] : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2177 = 5'h17 == rd ? _next_reg_T_65[31:0] : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2178 = 5'h18 == rd ? _next_reg_T_65[31:0] : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2179 = 5'h19 == rd ? _next_reg_T_65[31:0] : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2180 = 5'h1a == rd ? _next_reg_T_65[31:0] : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2181 = 5'h1b == rd ? _next_reg_T_65[31:0] : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2182 = 5'h1c == rd ? _next_reg_T_65[31:0] : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2183 = 5'h1d == rd ? _next_reg_T_65[31:0] : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2184 = 5'h1e == rd ? _next_reg_T_65[31:0] : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2185 = 5'h1f == rd ? _next_reg_T_65[31:0] : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _now_reg_rs1_35 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T_4 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 312:39]
  wire [31:0] _mem_read_addr_T_5 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 312:39]
  wire  _GEN_2186 = _T_437 | _GEN_2117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2187 = _T_437 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 312:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2188 = _T_437 ? 6'h20 : _GEN_2119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2189 = _T_437 ? _GEN_2154 : _GEN_2120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2190 = _T_437 ? _GEN_2155 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2191 = _T_437 ? _GEN_2156 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2192 = _T_437 ? _GEN_2157 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2193 = _T_437 ? _GEN_2158 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2194 = _T_437 ? _GEN_2159 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2195 = _T_437 ? _GEN_2160 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2196 = _T_437 ? _GEN_2161 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2197 = _T_437 ? _GEN_2162 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2198 = _T_437 ? _GEN_2163 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2199 = _T_437 ? _GEN_2164 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2200 = _T_437 ? _GEN_2165 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2201 = _T_437 ? _GEN_2166 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2202 = _T_437 ? _GEN_2167 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2203 = _T_437 ? _GEN_2168 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2204 = _T_437 ? _GEN_2169 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2205 = _T_437 ? _GEN_2170 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2206 = _T_437 ? _GEN_2171 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2207 = _T_437 ? _GEN_2172 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2208 = _T_437 ? _GEN_2173 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2209 = _T_437 ? _GEN_2174 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2210 = _T_437 ? _GEN_2175 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2211 = _T_437 ? _GEN_2176 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2212 = _T_437 ? _GEN_2177 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2213 = _T_437 ? _GEN_2178 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2214 = _T_437 ? _GEN_2179 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2215 = _T_437 ? _GEN_2180 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2216 = _T_437 ? _GEN_2181 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2217 = _T_437 ? _GEN_2182 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2218 = _T_437 ? _GEN_2183 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2219 = _T_437 ? _GEN_2184 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2220 = _T_437 ? _GEN_2185 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2222 = _T_437 ? _GEN_2153 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2226 = _T_388 ? inst[14:12] : _GEN_2113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2228 = _T_388 ? inst[6:0] : _GEN_2115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2230 = _T_388 ? _GEN_2186 : _GEN_2117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2231 = _T_388 ? _GEN_2187 : _GEN_2118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [5:0] _GEN_2232 = _T_388 ? _GEN_2188 : _GEN_2119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2233 = _T_388 ? _GEN_2189 : _GEN_2120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2234 = _T_388 ? _GEN_2190 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2235 = _T_388 ? _GEN_2191 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2236 = _T_388 ? _GEN_2192 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2237 = _T_388 ? _GEN_2193 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2238 = _T_388 ? _GEN_2194 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2239 = _T_388 ? _GEN_2195 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2240 = _T_388 ? _GEN_2196 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2241 = _T_388 ? _GEN_2197 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2242 = _T_388 ? _GEN_2198 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2243 = _T_388 ? _GEN_2199 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2244 = _T_388 ? _GEN_2200 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2245 = _T_388 ? _GEN_2201 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2246 = _T_388 ? _GEN_2202 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2247 = _T_388 ? _GEN_2203 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2248 = _T_388 ? _GEN_2204 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2249 = _T_388 ? _GEN_2205 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2250 = _T_388 ? _GEN_2206 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2251 = _T_388 ? _GEN_2207 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2252 = _T_388 ? _GEN_2208 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2253 = _T_388 ? _GEN_2209 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2254 = _T_388 ? _GEN_2210 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2255 = _T_388 ? _GEN_2211 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2256 = _T_388 ? _GEN_2212 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2257 = _T_388 ? _GEN_2213 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2258 = _T_388 ? _GEN_2214 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2259 = _T_388 ? _GEN_2215 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2260 = _T_388 ? _GEN_2216 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2261 = _T_388 ? _GEN_2217 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2262 = _T_388 ? _GEN_2218 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2263 = _T_388 ? _GEN_2219 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2264 = _T_388 ? _GEN_2220 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2266 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [2:0] _funct3_T_29 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_412 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _GEN_2268 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _now_reg_rs1_36 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_68 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:118]
  wire [31:0] _next_reg_T_69 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:118]
  wire [1:0] _next_reg_rOff_T_3 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_3 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_21 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_22 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_23 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_24 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_25 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_26 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_27 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_3 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_70 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6210 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_71 = _GEN_6207 & 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [7:0] _next_reg_T_72 = _next_reg_T_49[7:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:129]
  wire [31:0] _next_reg_T_73 = {24'h0,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_reg_rd_25 = {24'h0,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_2269 = 5'h0 == rd ? _next_reg_T_73 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2270 = 5'h1 == rd ? _next_reg_T_73 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2271 = 5'h2 == rd ? _next_reg_T_73 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2272 = 5'h3 == rd ? _next_reg_T_73 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2273 = 5'h4 == rd ? _next_reg_T_73 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2274 = 5'h5 == rd ? _next_reg_T_73 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2275 = 5'h6 == rd ? _next_reg_T_73 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2276 = 5'h7 == rd ? _next_reg_T_73 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2277 = 5'h8 == rd ? _next_reg_T_73 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2278 = 5'h9 == rd ? _next_reg_T_73 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2279 = 5'ha == rd ? _next_reg_T_73 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2280 = 5'hb == rd ? _next_reg_T_73 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2281 = 5'hc == rd ? _next_reg_T_73 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2282 = 5'hd == rd ? _next_reg_T_73 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2283 = 5'he == rd ? _next_reg_T_73 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2284 = 5'hf == rd ? _next_reg_T_73 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2285 = 5'h10 == rd ? _next_reg_T_73 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2286 = 5'h11 == rd ? _next_reg_T_73 : _GEN_2250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2287 = 5'h12 == rd ? _next_reg_T_73 : _GEN_2251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2288 = 5'h13 == rd ? _next_reg_T_73 : _GEN_2252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2289 = 5'h14 == rd ? _next_reg_T_73 : _GEN_2253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2290 = 5'h15 == rd ? _next_reg_T_73 : _GEN_2254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2291 = 5'h16 == rd ? _next_reg_T_73 : _GEN_2255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2292 = 5'h17 == rd ? _next_reg_T_73 : _GEN_2256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2293 = 5'h18 == rd ? _next_reg_T_73 : _GEN_2257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2294 = 5'h19 == rd ? _next_reg_T_73 : _GEN_2258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2295 = 5'h1a == rd ? _next_reg_T_73 : _GEN_2259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2296 = 5'h1b == rd ? _next_reg_T_73 : _GEN_2260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2297 = 5'h1c == rd ? _next_reg_T_73 : _GEN_2261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2298 = 5'h1d == rd ? _next_reg_T_73 : _GEN_2262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2299 = 5'h1e == rd ? _next_reg_T_73 : _GEN_2263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2300 = 5'h1f == rd ? _next_reg_T_73 : _GEN_2264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [2:0] _GEN_2304 = _T_408 ? inst[14:12] : _GEN_2226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2306 = _T_408 ? inst[6:0] : _GEN_2228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2309 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2310 = _T_408 | _GEN_2230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2311 = _T_408 ? _T_433 : _GEN_2231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2312 = _T_408 ? 6'h8 : _GEN_2232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2313 = _T_408 ? _GEN_2269 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2314 = _T_408 ? _GEN_2270 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2315 = _T_408 ? _GEN_2271 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2316 = _T_408 ? _GEN_2272 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2317 = _T_408 ? _GEN_2273 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2318 = _T_408 ? _GEN_2274 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2319 = _T_408 ? _GEN_2275 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2320 = _T_408 ? _GEN_2276 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2321 = _T_408 ? _GEN_2277 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2322 = _T_408 ? _GEN_2278 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2323 = _T_408 ? _GEN_2279 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2324 = _T_408 ? _GEN_2280 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2325 = _T_408 ? _GEN_2281 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2326 = _T_408 ? _GEN_2282 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2327 = _T_408 ? _GEN_2283 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2328 = _T_408 ? _GEN_2284 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2329 = _T_408 ? _GEN_2285 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2330 = _T_408 ? _GEN_2286 : _GEN_2250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2331 = _T_408 ? _GEN_2287 : _GEN_2251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2332 = _T_408 ? _GEN_2288 : _GEN_2252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2333 = _T_408 ? _GEN_2289 : _GEN_2253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2334 = _T_408 ? _GEN_2290 : _GEN_2254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2335 = _T_408 ? _GEN_2291 : _GEN_2255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2336 = _T_408 ? _GEN_2292 : _GEN_2256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2337 = _T_408 ? _GEN_2293 : _GEN_2257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2338 = _T_408 ? _GEN_2294 : _GEN_2258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2339 = _T_408 ? _GEN_2295 : _GEN_2259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2340 = _T_408 ? _GEN_2296 : _GEN_2260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2341 = _T_408 ? _GEN_2297 : _GEN_2261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2342 = _T_408 ? _GEN_2298 : _GEN_2262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2343 = _T_408 ? _GEN_2299 : _GEN_2263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2344 = _T_408 ? _GEN_2300 : _GEN_2264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [2:0] _funct3_T_30 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_431 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_38 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_74 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:54]
  wire [31:0] _next_reg_T_75 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:54]
  wire [1:0] _next_reg_rOff_T_4 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_4 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_28 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_29 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_30 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_31 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_32 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_33 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_34 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_4 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_76 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6211 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_77 = _GEN_6207 & 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [15:0] _next_reg_T_78 = _next_reg_T_57[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:66]
  wire [31:0] _next_reg_T_79 = {16'h0,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_reg_rd_26 = {16'h0,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_2345 = 5'h0 == rd ? _next_reg_T_79 : _GEN_2313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2346 = 5'h1 == rd ? _next_reg_T_79 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2347 = 5'h2 == rd ? _next_reg_T_79 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2348 = 5'h3 == rd ? _next_reg_T_79 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2349 = 5'h4 == rd ? _next_reg_T_79 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2350 = 5'h5 == rd ? _next_reg_T_79 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2351 = 5'h6 == rd ? _next_reg_T_79 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2352 = 5'h7 == rd ? _next_reg_T_79 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2353 = 5'h8 == rd ? _next_reg_T_79 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2354 = 5'h9 == rd ? _next_reg_T_79 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2355 = 5'ha == rd ? _next_reg_T_79 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2356 = 5'hb == rd ? _next_reg_T_79 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2357 = 5'hc == rd ? _next_reg_T_79 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2358 = 5'hd == rd ? _next_reg_T_79 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2359 = 5'he == rd ? _next_reg_T_79 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2360 = 5'hf == rd ? _next_reg_T_79 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2361 = 5'h10 == rd ? _next_reg_T_79 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2362 = 5'h11 == rd ? _next_reg_T_79 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2363 = 5'h12 == rd ? _next_reg_T_79 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2364 = 5'h13 == rd ? _next_reg_T_79 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2365 = 5'h14 == rd ? _next_reg_T_79 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2366 = 5'h15 == rd ? _next_reg_T_79 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2367 = 5'h16 == rd ? _next_reg_T_79 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2368 = 5'h17 == rd ? _next_reg_T_79 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2369 = 5'h18 == rd ? _next_reg_T_79 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2370 = 5'h19 == rd ? _next_reg_T_79 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2371 = 5'h1a == rd ? _next_reg_T_79 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2372 = 5'h1b == rd ? _next_reg_T_79 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2373 = 5'h1c == rd ? _next_reg_T_79 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2374 = 5'h1d == rd ? _next_reg_T_79 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2375 = 5'h1e == rd ? _next_reg_T_79 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2376 = 5'h1f == rd ? _next_reg_T_79 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _now_reg_rs1_39 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T_6 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 322:39]
  wire [31:0] _mem_read_addr_T_7 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 322:39]
  wire  _GEN_2377 = _T_435 | _GEN_2310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2378 = _T_435 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 322:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2379 = _T_435 ? 6'h10 : _GEN_2312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2380 = _T_435 ? _GEN_2345 : _GEN_2313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2381 = _T_435 ? _GEN_2346 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2382 = _T_435 ? _GEN_2347 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2383 = _T_435 ? _GEN_2348 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2384 = _T_435 ? _GEN_2349 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2385 = _T_435 ? _GEN_2350 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2386 = _T_435 ? _GEN_2351 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2387 = _T_435 ? _GEN_2352 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2388 = _T_435 ? _GEN_2353 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2389 = _T_435 ? _GEN_2354 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2390 = _T_435 ? _GEN_2355 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2391 = _T_435 ? _GEN_2356 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2392 = _T_435 ? _GEN_2357 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2393 = _T_435 ? _GEN_2358 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2394 = _T_435 ? _GEN_2359 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2395 = _T_435 ? _GEN_2360 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2396 = _T_435 ? _GEN_2361 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2397 = _T_435 ? _GEN_2362 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2398 = _T_435 ? _GEN_2363 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2399 = _T_435 ? _GEN_2364 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2400 = _T_435 ? _GEN_2365 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2401 = _T_435 ? _GEN_2366 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2402 = _T_435 ? _GEN_2367 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2403 = _T_435 ? _GEN_2368 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2404 = _T_435 ? _GEN_2369 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2405 = _T_435 ? _GEN_2370 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2406 = _T_435 ? _GEN_2371 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2407 = _T_435 ? _GEN_2372 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2408 = _T_435 ? _GEN_2373 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2409 = _T_435 ? _GEN_2374 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2410 = _T_435 ? _GEN_2375 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2411 = _T_435 ? _GEN_2376 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_2413 = _T_435 ? _GEN_2266 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2417 = _T_427 ? inst[14:12] : _GEN_2304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2419 = _T_427 ? inst[6:0] : _GEN_2306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2421 = _T_427 ? _GEN_2377 : _GEN_2310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2422 = _T_427 ? _GEN_2074 : _GEN_2311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [5:0] _GEN_2423 = _T_427 ? _GEN_2379 : _GEN_2312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2424 = _T_427 ? _GEN_2380 : _GEN_2313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2425 = _T_427 ? _GEN_2381 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2426 = _T_427 ? _GEN_2382 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2427 = _T_427 ? _GEN_2383 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2428 = _T_427 ? _GEN_2384 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2429 = _T_427 ? _GEN_2385 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2430 = _T_427 ? _GEN_2386 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2431 = _T_427 ? _GEN_2387 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2432 = _T_427 ? _GEN_2388 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2433 = _T_427 ? _GEN_2389 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2434 = _T_427 ? _GEN_2390 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2435 = _T_427 ? _GEN_2391 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2436 = _T_427 ? _GEN_2392 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2437 = _T_427 ? _GEN_2393 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2438 = _T_427 ? _GEN_2394 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2439 = _T_427 ? _GEN_2395 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2440 = _T_427 ? _GEN_2396 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2441 = _T_427 ? _GEN_2397 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2442 = _T_427 ? _GEN_2398 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2443 = _T_427 ? _GEN_2399 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2444 = _T_427 ? _GEN_2400 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2445 = _T_427 ? _GEN_2401 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2446 = _T_427 ? _GEN_2402 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2447 = _T_427 ? _GEN_2403 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2448 = _T_427 ? _GEN_2404 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2449 = _T_427 ? _GEN_2405 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2450 = _T_427 ? _GEN_2406 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2451 = _T_427 ? _GEN_2407 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2452 = _T_427 ? _GEN_2408 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2453 = _T_427 ? _GEN_2409 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2454 = _T_427 ? _GEN_2410 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2455 = _T_427 ? _GEN_2411 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_2457 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [2:0] _funct3_T_31 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_452 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _GEN_2459 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _now_reg_rs1_40 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_466 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:95]
  wire [31:0] _T_467 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:95]
  wire [31:0] _now_reg_rs2_15 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [7:0] _T_468 = _GEN_840[7:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:119]
  wire [2:0] _GEN_2464 = _T_447 ? inst[14:12] : _GEN_2417; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2466 = _T_447 ? inst[6:0] : _GEN_2419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2469 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _mem_WIRE_write_valid = 1'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire  _GEN_2470 = 32'h23 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _mem_WIRE_write_addr = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [31:0] _GEN_2471 = _T_447 ? _T_433 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [5:0] _mem_WIRE_write_memWidth = 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [5:0] _GEN_2472 = _T_447 ? 6'h8 : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _mem_WIRE_write_data = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [31:0] _GEN_2473 = _T_447 ? {{24'd0}, _GEN_840[7:0]} : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [2:0] _funct3_T_32 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_475 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_42 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_490 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 331:31]
  wire [31:0] _T_491 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 331:31]
  wire [31:0] _now_reg_rs2_16 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [15:0] _T_492 = _GEN_840[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 331:56]
  wire [31:0] _now_reg_rs1_43 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_write_addr_T = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 333:40]
  wire [31:0] _mem_write_addr_T_1 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 333:40]
  wire  _GEN_2474 = _T_435 | _T_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [31:0] _GEN_2475 = _T_435 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 333:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [5:0] _GEN_2476 = _T_435 ? 6'h10 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [31:0] _GEN_2477 = _T_435 ? {{16'd0}, _GEN_840[15:0]} : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_2479 = _T_435 ? _GEN_2457 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2484 = _T_470 ? inst[14:12] : _GEN_2464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2486 = _T_470 ? inst[6:0] : _GEN_2466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2488 = _T_470 ? _GEN_2474 : _T_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [31:0] _GEN_2489 = _T_470 ? _GEN_2074 : _GEN_2471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [5:0] _GEN_2490 = _T_470 ? _GEN_2476 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [31:0] _GEN_2491 = _T_470 ? _GEN_2477 : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2493 = _T_470 ? _GEN_2479 : _GEN_2457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [2:0] _funct3_T_33 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_499 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_45 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_514 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 340:31]
  wire [31:0] _T_515 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 340:31]
  wire [31:0] _now_reg_rs2_17 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_516 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _now_reg_rs1_46 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_write_addr_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 342:40]
  wire [31:0] _mem_write_addr_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 342:40]
  wire  _GEN_2494 = _T_437 | _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [31:0] _GEN_2495 = _T_437 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 342:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [5:0] _GEN_2496 = _T_437 ? 6'h20 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [31:0] _GEN_2497 = _T_437 ? _GEN_840 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_2499 = _T_437 ? _GEN_2493 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2504 = _T_494 ? inst[14:12] : _GEN_2484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2506 = _T_494 ? inst[6:0] : _GEN_2486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2508 = _T_494 ? _GEN_2494 : _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [31:0] _GEN_2509 = _T_494 ? _GEN_2187 : _GEN_2489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [5:0] _GEN_2510 = _T_494 ? _GEN_2496 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [31:0] _GEN_2511 = _T_494 ? _GEN_2497 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_2513 = _T_494 ? _GEN_2499 : _GEN_2493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [2:0] _funct3_T_34 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_522 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_2517 = _T_518 ? inst[14:12] : _GEN_2504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2519 = _T_518 ? inst[6:0] : _GEN_2506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2522 = _T_518 | _GEN_2513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _funct3_T_35 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_528 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _GEN_2524 = 2'h0 == io_now_internal_privilegeMode | _GEN_2522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2526 = 2'h1 == io_now_internal_privilegeMode | (2'h0 == io_now_internal_privilegeMode | _GEN_2522); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2529 = 2'h3 == io_now_internal_privilegeMode | (2'h1 == io_now_internal_privilegeMode | (2'h0 ==
    io_now_internal_privilegeMode | _GEN_2522)); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2535 = _T_524 ? inst[14:12] : _GEN_2517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2537 = _T_524 ? inst[6:0] : _GEN_2519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2540 = _T_524 ? _GEN_2529 : _GEN_2522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23]
  wire [2:0] _funct3_T_36 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_537 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_2546 = _T_533 ? inst[14:12] : _GEN_2535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2548 = _T_533 ? inst[6:0] : _GEN_2537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [2:0] _funct3_T_37 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_546 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_547 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_reg_T_80 = io_now_reg_2 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:52]
  wire [31:0] _next_reg_T_81 = io_now_reg_2 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:52]
  wire [1:0] _next_reg_rOff_T_5 = _next_reg_T_81[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_5 = {_next_reg_T_81[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_35 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_36 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_37 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_38 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_39 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_40 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_41 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_5 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_82 = io_mem_read_data >> next_reg_rOff_5; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6212 = {{32'd0}, _next_reg_T_82}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_83 = _GEN_6212 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [31:0] _next_reg_T_84 = _next_reg_T_83[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:64]
  wire  next_reg_signBit_3 = _next_reg_T_83[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_85 = _next_reg_T_83[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:64]
  wire [31:0] _next_reg_rd_27 = _next_reg_T_83[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:64]
  wire [31:0] _GEN_2550 = 5'h0 == rd ? _next_reg_T_83[31:0] : _GEN_2424; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2551 = 5'h1 == rd ? _next_reg_T_83[31:0] : _GEN_2425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2552 = 5'h2 == rd ? _next_reg_T_83[31:0] : _GEN_2426; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2553 = 5'h3 == rd ? _next_reg_T_83[31:0] : _GEN_2427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2554 = 5'h4 == rd ? _next_reg_T_83[31:0] : _GEN_2428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2555 = 5'h5 == rd ? _next_reg_T_83[31:0] : _GEN_2429; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2556 = 5'h6 == rd ? _next_reg_T_83[31:0] : _GEN_2430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2557 = 5'h7 == rd ? _next_reg_T_83[31:0] : _GEN_2431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2558 = 5'h8 == rd ? _next_reg_T_83[31:0] : _GEN_2432; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2559 = 5'h9 == rd ? _next_reg_T_83[31:0] : _GEN_2433; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2560 = 5'ha == rd ? _next_reg_T_83[31:0] : _GEN_2434; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2561 = 5'hb == rd ? _next_reg_T_83[31:0] : _GEN_2435; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2562 = 5'hc == rd ? _next_reg_T_83[31:0] : _GEN_2436; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2563 = 5'hd == rd ? _next_reg_T_83[31:0] : _GEN_2437; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2564 = 5'he == rd ? _next_reg_T_83[31:0] : _GEN_2438; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2565 = 5'hf == rd ? _next_reg_T_83[31:0] : _GEN_2439; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2566 = 5'h10 == rd ? _next_reg_T_83[31:0] : _GEN_2440; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2567 = 5'h11 == rd ? _next_reg_T_83[31:0] : _GEN_2441; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2568 = 5'h12 == rd ? _next_reg_T_83[31:0] : _GEN_2442; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2569 = 5'h13 == rd ? _next_reg_T_83[31:0] : _GEN_2443; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2570 = 5'h14 == rd ? _next_reg_T_83[31:0] : _GEN_2444; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2571 = 5'h15 == rd ? _next_reg_T_83[31:0] : _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2572 = 5'h16 == rd ? _next_reg_T_83[31:0] : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2573 = 5'h17 == rd ? _next_reg_T_83[31:0] : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2574 = 5'h18 == rd ? _next_reg_T_83[31:0] : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2575 = 5'h19 == rd ? _next_reg_T_83[31:0] : _GEN_2449; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2576 = 5'h1a == rd ? _next_reg_T_83[31:0] : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2577 = 5'h1b == rd ? _next_reg_T_83[31:0] : _GEN_2451; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2578 = 5'h1c == rd ? _next_reg_T_83[31:0] : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2579 = 5'h1d == rd ? _next_reg_T_83[31:0] : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2580 = 5'h1e == rd ? _next_reg_T_83[31:0] : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [31:0] _GEN_2581 = 5'h1f == rd ? _next_reg_T_83[31:0] : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [2:0] _GEN_2583 = _T_542 ? inst[15:13] : _GEN_2546; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_2584 = _T_542 & inst[12]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:22]
  wire [4:0] _GEN_2586 = _T_542 ? inst[6:2] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:52]
  wire [1:0] _GEN_2587 = _T_542 ? inst[1:0] : 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 97:24]
  wire  _GEN_2590 = _T_542 | _GEN_2421; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2591 = _T_542 ? _next_reg_T_81 : _GEN_2422; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2592 = _T_542 ? 6'h20 : _GEN_2423; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2593 = _T_542 ? _GEN_2550 : _GEN_2424; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2594 = _T_542 ? _GEN_2551 : _GEN_2425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2595 = _T_542 ? _GEN_2552 : _GEN_2426; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2596 = _T_542 ? _GEN_2553 : _GEN_2427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2597 = _T_542 ? _GEN_2554 : _GEN_2428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2598 = _T_542 ? _GEN_2555 : _GEN_2429; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2599 = _T_542 ? _GEN_2556 : _GEN_2430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2600 = _T_542 ? _GEN_2557 : _GEN_2431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2601 = _T_542 ? _GEN_2558 : _GEN_2432; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2602 = _T_542 ? _GEN_2559 : _GEN_2433; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2603 = _T_542 ? _GEN_2560 : _GEN_2434; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2604 = _T_542 ? _GEN_2561 : _GEN_2435; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2605 = _T_542 ? _GEN_2562 : _GEN_2436; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2606 = _T_542 ? _GEN_2563 : _GEN_2437; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2607 = _T_542 ? _GEN_2564 : _GEN_2438; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2608 = _T_542 ? _GEN_2565 : _GEN_2439; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2609 = _T_542 ? _GEN_2566 : _GEN_2440; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2610 = _T_542 ? _GEN_2567 : _GEN_2441; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2611 = _T_542 ? _GEN_2568 : _GEN_2442; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2612 = _T_542 ? _GEN_2569 : _GEN_2443; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2613 = _T_542 ? _GEN_2570 : _GEN_2444; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2614 = _T_542 ? _GEN_2571 : _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2615 = _T_542 ? _GEN_2572 : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2616 = _T_542 ? _GEN_2573 : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2617 = _T_542 ? _GEN_2574 : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2618 = _T_542 ? _GEN_2575 : _GEN_2449; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2619 = _T_542 ? _GEN_2576 : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2620 = _T_542 ? _GEN_2577 : _GEN_2451; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2621 = _T_542 ? _GEN_2578 : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2622 = _T_542 ? _GEN_2579 : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2623 = _T_542 ? _GEN_2580 : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [31:0] _GEN_2624 = _T_542 ? _GEN_2581 : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [2:0] _funct3_T_38 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _ph6_T = inst[12:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_553 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _T_554 = io_now_reg_2 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 146:29]
  wire [31:0] _T_555 = io_now_reg_2 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 146:29]
  wire [31:0] _now_reg_rs2_18 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_556 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [2:0] _GEN_2626 = _T_549 ? inst[15:13] : _GEN_2583; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_2627 = _T_549 ? inst[12:7] : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 104:22]
  wire [1:0] _GEN_2629 = _T_549 ? inst[1:0] : _GEN_2587; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2631 = _T_549 | _GEN_2508; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [31:0] _GEN_2632 = _T_549 ? _next_reg_T_81 : _GEN_2509; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [5:0] _GEN_2633 = _T_549 ? 6'h20 : _GEN_2510; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [31:0] _GEN_2634 = _T_549 ? _GEN_840 : _GEN_2511; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire [15:0] _T_559 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 116:97]
  wire [2:0] _funct3_T_39 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [12:0] _T_560 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _ph3_T = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [9:0] _T_561 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_562 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [1:0] _ph2_T = inst[6:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _T_563 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rdP_T = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_564 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [15:0] _T_798 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:97]
  wire [9:0] _T_799 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_10 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_790 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:97]
  wire [9:0] _T_791 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_9 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_782 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:97]
  wire [9:0] _T_783 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_8 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_774 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:97]
  wire [9:0] _T_775 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_7 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_742 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:97]
  wire [12:0] _T_743 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [9:0] _T_744 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_6 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_734 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:97]
  wire [12:0] _T_735 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [9:0] _T_736 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_5 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_718 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:97]
  wire [12:0] _T_719 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [9:0] _T_720 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_4 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_618 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:97]
  wire [12:0] _T_619 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [9:0] _T_620 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_3 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_609 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:97]
  wire [12:0] _T_610 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [9:0] _T_611 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_2 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [15:0] _T_568 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 117:97]
  wire [12:0] _T_569 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [9:0] _T_570 = inst[9:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs1P_T_1 = inst[9:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _GEN_2702 = _T_558 ? inst[9:7] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [2:0] _GEN_2809 = _T_567 ? inst[9:7] : _GEN_2702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2887 = _T_608 ? inst[9:7] : _GEN_2809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2931 = _T_617 ? inst[9:7] : _GEN_2887; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3400 = _T_717 ? inst[9:7] : _GEN_2931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3504 = _T_733 ? inst[9:7] : _GEN_3400; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3608 = _T_741 ? inst[9:7] : _GEN_3504; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3883 = _T_773 ? inst[9:7] : _GEN_3608; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4018 = _T_781 ? inst[9:7] : _GEN_3883; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4153 = _T_789 ? inst[9:7] : _GEN_4018; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4288 = _T_797 ? inst[9:7] : _GEN_4153; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] rs1P = io_valid ? _GEN_4288 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [2:0] _GEN_6178 = rs1P; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [15:0] _T_685 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 115:97]
  wire [12:0] _T_686 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_687 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rdP_T_1 = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _GEN_2704 = _T_558 ? inst[4:2] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [2:0] _GEN_2890 = _T_608 ? rs1P : _GEN_2704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 186:24]
  wire [2:0] _GEN_2934 = _T_617 ? rs1P : _GEN_2890; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 194:24]
  wire [2:0] _GEN_3227 = _T_684 ? inst[4:2] : _GEN_2934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3403 = _T_717 ? rs1P : _GEN_3227; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 235:24]
  wire [2:0] _GEN_3507 = _T_733 ? rs1P : _GEN_3403; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 240:24]
  wire [2:0] _GEN_3611 = _T_741 ? rs1P : _GEN_3507; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 245:24]
  wire [2:0] _GEN_3887 = _T_773 ? rs1P : _GEN_3611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 253:23]
  wire [2:0] _GEN_4022 = _T_781 ? rs1P : _GEN_3887; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 254:23]
  wire [2:0] _GEN_4157 = _T_789 ? rs1P : _GEN_4022; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 255:23]
  wire [2:0] _GEN_4292 = _T_797 ? rs1P : _GEN_4157; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 256:23]
  wire [2:0] rdP = io_valid ? _GEN_4292 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [2:0] _GEN_6180 = rdP; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [4:0] _T_565 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_86 = {2'h1,rs1P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_2635 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_2636 = 5'h1 == _next_reg_T_86 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2637 = 5'h2 == _next_reg_T_86 ? io_now_reg_2 : _GEN_2636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2638 = 5'h3 == _next_reg_T_86 ? io_now_reg_3 : _GEN_2637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2639 = 5'h4 == _next_reg_T_86 ? io_now_reg_4 : _GEN_2638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2640 = 5'h5 == _next_reg_T_86 ? io_now_reg_5 : _GEN_2639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2641 = 5'h6 == _next_reg_T_86 ? io_now_reg_6 : _GEN_2640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2642 = 5'h7 == _next_reg_T_86 ? io_now_reg_7 : _GEN_2641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2643 = 5'h8 == _next_reg_T_86 ? io_now_reg_8 : _GEN_2642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2644 = 5'h9 == _next_reg_T_86 ? io_now_reg_9 : _GEN_2643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2645 = 5'ha == _next_reg_T_86 ? io_now_reg_10 : _GEN_2644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2646 = 5'hb == _next_reg_T_86 ? io_now_reg_11 : _GEN_2645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2647 = 5'hc == _next_reg_T_86 ? io_now_reg_12 : _GEN_2646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2648 = 5'hd == _next_reg_T_86 ? io_now_reg_13 : _GEN_2647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2649 = 5'he == _next_reg_T_86 ? io_now_reg_14 : _GEN_2648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2650 = 5'hf == _next_reg_T_86 ? io_now_reg_15 : _GEN_2649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2651 = 5'h10 == _next_reg_T_86 ? io_now_reg_16 : _GEN_2650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2652 = 5'h11 == _next_reg_T_86 ? io_now_reg_17 : _GEN_2651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2653 = 5'h12 == _next_reg_T_86 ? io_now_reg_18 : _GEN_2652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2654 = 5'h13 == _next_reg_T_86 ? io_now_reg_19 : _GEN_2653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2655 = 5'h14 == _next_reg_T_86 ? io_now_reg_20 : _GEN_2654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2656 = 5'h15 == _next_reg_T_86 ? io_now_reg_21 : _GEN_2655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2657 = 5'h16 == _next_reg_T_86 ? io_now_reg_22 : _GEN_2656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2658 = 5'h17 == _next_reg_T_86 ? io_now_reg_23 : _GEN_2657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2659 = 5'h18 == _next_reg_T_86 ? io_now_reg_24 : _GEN_2658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2660 = 5'h19 == _next_reg_T_86 ? io_now_reg_25 : _GEN_2659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2661 = 5'h1a == _next_reg_T_86 ? io_now_reg_26 : _GEN_2660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2662 = 5'h1b == _next_reg_T_86 ? io_now_reg_27 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2663 = 5'h1c == _next_reg_T_86 ? io_now_reg_28 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2664 = 5'h1d == _next_reg_T_86 ? io_now_reg_29 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2665 = 5'h1e == _next_reg_T_86 ? io_now_reg_30 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _GEN_2666 = 5'h1f == _next_reg_T_86 ? io_now_reg_31 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [31:0] _now_reg_next_reg_T_86 = 5'h1f == _next_reg_T_86 ? io_now_reg_31 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [32:0] _next_reg_T_87 = _GEN_2666 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:68]
  wire [31:0] _next_reg_T_88 = _GEN_2666 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:68]
  wire [1:0] _next_reg_rOff_T_6 = _next_reg_T_88[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_6 = {_next_reg_T_88[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_42 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_43 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_44 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_45 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_46 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_47 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_48 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_6 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_89 = io_mem_read_data >> next_reg_rOff_6; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_6213 = {{32'd0}, _next_reg_T_89}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_90 = _GEN_6213 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [31:0] _next_reg_T_91 = _next_reg_T_90[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:80]
  wire  next_reg_signBit_4 = _next_reg_T_90[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_92 = _next_reg_T_90[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:80]
  wire [31:0] _next_reg_T_565 = _next_reg_T_90[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:80]
  wire [31:0] _GEN_2667 = 5'h0 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2593; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2668 = 5'h1 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2594; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2669 = 5'h2 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2595; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2670 = 5'h3 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2596; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2671 = 5'h4 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2597; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2672 = 5'h5 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2598; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2673 = 5'h6 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2599; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2674 = 5'h7 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2600; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2675 = 5'h8 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2601; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2676 = 5'h9 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2602; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2677 = 5'ha == _T_565 ? _next_reg_T_90[31:0] : _GEN_2603; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2678 = 5'hb == _T_565 ? _next_reg_T_90[31:0] : _GEN_2604; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2679 = 5'hc == _T_565 ? _next_reg_T_90[31:0] : _GEN_2605; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2680 = 5'hd == _T_565 ? _next_reg_T_90[31:0] : _GEN_2606; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2681 = 5'he == _T_565 ? _next_reg_T_90[31:0] : _GEN_2607; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2682 = 5'hf == _T_565 ? _next_reg_T_90[31:0] : _GEN_2608; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2683 = 5'h10 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2609; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2684 = 5'h11 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2685 = 5'h12 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2686 = 5'h13 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2612; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2687 = 5'h14 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2688 = 5'h15 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2689 = 5'h16 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2690 = 5'h17 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2691 = 5'h18 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2692 = 5'h19 == _T_565 ? _next_reg_T_90[31:0] : _GEN_2618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2693 = 5'h1a == _T_565 ? _next_reg_T_90[31:0] : _GEN_2619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2694 = 5'h1b == _T_565 ? _next_reg_T_90[31:0] : _GEN_2620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2695 = 5'h1c == _T_565 ? _next_reg_T_90[31:0] : _GEN_2621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2696 = 5'h1d == _T_565 ? _next_reg_T_90[31:0] : _GEN_2622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2697 = 5'h1e == _T_565 ? _next_reg_T_90[31:0] : _GEN_2623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [31:0] _GEN_2698 = 5'h1f == _T_565 ? _next_reg_T_90[31:0] : _GEN_2624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [2:0] _GEN_2700 = _T_558 ? inst[15:13] : _GEN_2626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2701 = _T_558 ? inst[12:10] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:22]
  wire [1:0] _GEN_2703 = _T_558 ? inst[6:5] : 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:52]
  wire [1:0] _GEN_2705 = _T_558 ? inst[1:0] : _GEN_2629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2707 = _T_558 | _GEN_2590; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2708 = _T_558 ? _next_reg_T_88 : _GEN_2591; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2709 = _T_558 ? 6'h20 : _GEN_2592; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2710 = _T_558 ? _GEN_2667 : _GEN_2593; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2711 = _T_558 ? _GEN_2668 : _GEN_2594; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2712 = _T_558 ? _GEN_2669 : _GEN_2595; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2713 = _T_558 ? _GEN_2670 : _GEN_2596; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2714 = _T_558 ? _GEN_2671 : _GEN_2597; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2715 = _T_558 ? _GEN_2672 : _GEN_2598; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2716 = _T_558 ? _GEN_2673 : _GEN_2599; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2717 = _T_558 ? _GEN_2674 : _GEN_2600; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2718 = _T_558 ? _GEN_2675 : _GEN_2601; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2719 = _T_558 ? _GEN_2676 : _GEN_2602; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2720 = _T_558 ? _GEN_2677 : _GEN_2603; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2721 = _T_558 ? _GEN_2678 : _GEN_2604; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2722 = _T_558 ? _GEN_2679 : _GEN_2605; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2723 = _T_558 ? _GEN_2680 : _GEN_2606; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2724 = _T_558 ? _GEN_2681 : _GEN_2607; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2725 = _T_558 ? _GEN_2682 : _GEN_2608; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2726 = _T_558 ? _GEN_2683 : _GEN_2609; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2727 = _T_558 ? _GEN_2684 : _GEN_2610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2728 = _T_558 ? _GEN_2685 : _GEN_2611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2729 = _T_558 ? _GEN_2686 : _GEN_2612; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2730 = _T_558 ? _GEN_2687 : _GEN_2613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2731 = _T_558 ? _GEN_2688 : _GEN_2614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2732 = _T_558 ? _GEN_2689 : _GEN_2615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2733 = _T_558 ? _GEN_2690 : _GEN_2616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2734 = _T_558 ? _GEN_2691 : _GEN_2617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2735 = _T_558 ? _GEN_2692 : _GEN_2618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2736 = _T_558 ? _GEN_2693 : _GEN_2619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2737 = _T_558 ? _GEN_2694 : _GEN_2620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2738 = _T_558 ? _GEN_2695 : _GEN_2621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2739 = _T_558 ? _GEN_2696 : _GEN_2622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2740 = _T_558 ? _GEN_2697 : _GEN_2623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [31:0] _GEN_2741 = _T_558 ? _GEN_2698 : _GEN_2624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [2:0] _funct3_T_40 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _ph3_T_1 = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_571 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [1:0] _ph2_T_1 = inst[6:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _T_572 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs2P_T = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_573 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_574 = {2'h1,rs1P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_2742 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_2743 = 5'h1 == _next_reg_T_86 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2744 = 5'h2 == _next_reg_T_86 ? io_now_reg_2 : _GEN_2636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2745 = 5'h3 == _next_reg_T_86 ? io_now_reg_3 : _GEN_2637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2746 = 5'h4 == _next_reg_T_86 ? io_now_reg_4 : _GEN_2638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2747 = 5'h5 == _next_reg_T_86 ? io_now_reg_5 : _GEN_2639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2748 = 5'h6 == _next_reg_T_86 ? io_now_reg_6 : _GEN_2640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2749 = 5'h7 == _next_reg_T_86 ? io_now_reg_7 : _GEN_2641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2750 = 5'h8 == _next_reg_T_86 ? io_now_reg_8 : _GEN_2642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2751 = 5'h9 == _next_reg_T_86 ? io_now_reg_9 : _GEN_2643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2752 = 5'ha == _next_reg_T_86 ? io_now_reg_10 : _GEN_2644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2753 = 5'hb == _next_reg_T_86 ? io_now_reg_11 : _GEN_2645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2754 = 5'hc == _next_reg_T_86 ? io_now_reg_12 : _GEN_2646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2755 = 5'hd == _next_reg_T_86 ? io_now_reg_13 : _GEN_2647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2756 = 5'he == _next_reg_T_86 ? io_now_reg_14 : _GEN_2648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2757 = 5'hf == _next_reg_T_86 ? io_now_reg_15 : _GEN_2649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2758 = 5'h10 == _next_reg_T_86 ? io_now_reg_16 : _GEN_2650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2759 = 5'h11 == _next_reg_T_86 ? io_now_reg_17 : _GEN_2651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2760 = 5'h12 == _next_reg_T_86 ? io_now_reg_18 : _GEN_2652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2761 = 5'h13 == _next_reg_T_86 ? io_now_reg_19 : _GEN_2653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2762 = 5'h14 == _next_reg_T_86 ? io_now_reg_20 : _GEN_2654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2763 = 5'h15 == _next_reg_T_86 ? io_now_reg_21 : _GEN_2655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2764 = 5'h16 == _next_reg_T_86 ? io_now_reg_22 : _GEN_2656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2765 = 5'h17 == _next_reg_T_86 ? io_now_reg_23 : _GEN_2657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2766 = 5'h18 == _next_reg_T_86 ? io_now_reg_24 : _GEN_2658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2767 = 5'h19 == _next_reg_T_86 ? io_now_reg_25 : _GEN_2659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2768 = 5'h1a == _next_reg_T_86 ? io_now_reg_26 : _GEN_2660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2769 = 5'h1b == _next_reg_T_86 ? io_now_reg_27 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2770 = 5'h1c == _next_reg_T_86 ? io_now_reg_28 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2771 = 5'h1d == _next_reg_T_86 ? io_now_reg_29 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2772 = 5'h1e == _next_reg_T_86 ? io_now_reg_30 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _GEN_2773 = 5'h1f == _next_reg_T_86 ? io_now_reg_31 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [31:0] _now_reg_T_574 = _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:{37,37}]
  wire [32:0] _T_575 = _GEN_2666 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:37]
  wire [31:0] _T_576 = _GEN_2666 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 157:37]
  wire [6:0] _T_800 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_801 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs2P_T_4 = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_792 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_793 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs2P_T_3 = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_784 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_785 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs2P_T_2 = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_776 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_777 = inst[4:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _rs2P_T_1 = inst[4:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _GEN_2811 = _T_567 ? inst[4:2] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [2:0] _GEN_3885 = _T_773 ? inst[4:2] : _GEN_2811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4020 = _T_781 ? inst[4:2] : _GEN_3885; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4155 = _T_789 ? inst[4:2] : _GEN_4020; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4290 = _T_797 ? inst[4:2] : _GEN_4155; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] rs2P = io_valid ? _GEN_4290 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [2:0] _GEN_6181 = rs2P; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [4:0] _T_577 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_2774 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_2775 = 5'h1 == _T_577 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2776 = 5'h2 == _T_577 ? io_now_reg_2 : _GEN_2775; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2777 = 5'h3 == _T_577 ? io_now_reg_3 : _GEN_2776; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2778 = 5'h4 == _T_577 ? io_now_reg_4 : _GEN_2777; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2779 = 5'h5 == _T_577 ? io_now_reg_5 : _GEN_2778; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2780 = 5'h6 == _T_577 ? io_now_reg_6 : _GEN_2779; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2781 = 5'h7 == _T_577 ? io_now_reg_7 : _GEN_2780; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2782 = 5'h8 == _T_577 ? io_now_reg_8 : _GEN_2781; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2783 = 5'h9 == _T_577 ? io_now_reg_9 : _GEN_2782; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2784 = 5'ha == _T_577 ? io_now_reg_10 : _GEN_2783; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2785 = 5'hb == _T_577 ? io_now_reg_11 : _GEN_2784; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2786 = 5'hc == _T_577 ? io_now_reg_12 : _GEN_2785; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2787 = 5'hd == _T_577 ? io_now_reg_13 : _GEN_2786; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2788 = 5'he == _T_577 ? io_now_reg_14 : _GEN_2787; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2789 = 5'hf == _T_577 ? io_now_reg_15 : _GEN_2788; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2790 = 5'h10 == _T_577 ? io_now_reg_16 : _GEN_2789; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2791 = 5'h11 == _T_577 ? io_now_reg_17 : _GEN_2790; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2792 = 5'h12 == _T_577 ? io_now_reg_18 : _GEN_2791; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2793 = 5'h13 == _T_577 ? io_now_reg_19 : _GEN_2792; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2794 = 5'h14 == _T_577 ? io_now_reg_20 : _GEN_2793; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2795 = 5'h15 == _T_577 ? io_now_reg_21 : _GEN_2794; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2796 = 5'h16 == _T_577 ? io_now_reg_22 : _GEN_2795; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2797 = 5'h17 == _T_577 ? io_now_reg_23 : _GEN_2796; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2798 = 5'h18 == _T_577 ? io_now_reg_24 : _GEN_2797; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2799 = 5'h19 == _T_577 ? io_now_reg_25 : _GEN_2798; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2800 = 5'h1a == _T_577 ? io_now_reg_26 : _GEN_2799; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2801 = 5'h1b == _T_577 ? io_now_reg_27 : _GEN_2800; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2802 = 5'h1c == _T_577 ? io_now_reg_28 : _GEN_2801; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2803 = 5'h1d == _T_577 ? io_now_reg_29 : _GEN_2802; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2804 = 5'h1e == _T_577 ? io_now_reg_30 : _GEN_2803; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2805 = 5'h1f == _T_577 ? io_now_reg_31 : _GEN_2804; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [2:0] _GEN_2807 = _T_567 ? inst[15:13] : _GEN_2700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2808 = _T_567 ? inst[12:10] : _GEN_2701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2810 = _T_567 ? inst[6:5] : _GEN_2703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2812 = _T_567 ? inst[1:0] : _GEN_2705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2814 = _T_567 | _GEN_2631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [31:0] _GEN_2815 = _T_567 ? _next_reg_T_88 : _GEN_2632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [5:0] _GEN_2816 = _T_567 ? 6'h20 : _GEN_2633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [31:0] _now_reg_T_577 = 5'h1f == _T_577 ? io_now_reg_31 : _GEN_2804; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [31:0] _GEN_2817 = _T_567 ? _GEN_2805 : _GEN_2634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire [15:0] _T_580 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 120:97]
  wire [2:0] _funct3_T_41 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [12:0] _T_581 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [10:0] _ph11_T = inst[12:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_582 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_18 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 164:35]
  wire [31:0] _next_pc_T_19 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 164:35]
  wire [2:0] _GEN_2819 = _T_579 ? inst[15:13] : _GEN_2807; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [10:0] _GEN_2820 = _T_579 ? inst[12:2] : 11'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 107:22]
  wire [1:0] _GEN_2821 = _T_579 ? inst[1:0] : _GEN_2812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2823 = _T_579 | _GEN_1923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 163:25]
  wire [31:0] _GEN_2824 = _T_579 ? _T_334 : _GEN_1924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 164:25]
  wire [15:0] _T_586 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 120:97]
  wire [2:0] _funct3_T_42 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [12:0] _T_587 = inst[12:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [10:0] _ph11_T_1 = inst[12:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_588 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_20 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 170:35]
  wire [31:0] _next_pc_T_21 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 170:35]
  wire [32:0] _next_reg_1_T = io_now_pc + 32'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 171:35]
  wire [31:0] _next_reg_1_T_1 = io_now_pc + 32'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 171:35]
  wire [2:0] _GEN_2826 = _T_584 ? inst[15:13] : _GEN_2819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [10:0] _GEN_2827 = _T_584 ? inst[12:2] : _GEN_2820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2828 = _T_584 ? inst[1:0] : _GEN_2821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2830 = _T_584 | _GEN_2823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 169:25]
  wire [31:0] _GEN_2831 = _T_584 ? _T_334 : _GEN_2824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 170:25]
  wire [31:0] _GEN_2832 = _T_584 ? _next_reg_1_T_1 : _GEN_2711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 166:23 171:25]
  wire [3:0] _funct4_T = inst[15:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_597 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_47 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [30:0] _next_pc_T_22 = _GEN_31[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 177:34]
  wire [31:0] _next_pc_T_23 = {_GEN_31[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 177:21]
  wire [3:0] _GEN_2834 = _T_593 ? inst[15:12] : 4'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 95:24]
  wire [1:0] _GEN_2837 = _T_593 ? inst[1:0] : _GEN_2828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2839 = _T_593 | _GEN_2830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 175:25]
  wire [31:0] _GEN_2840 = _T_593 ? _next_pc_T_23 : _GEN_2831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 177:15]
  wire [3:0] _funct4_T_1 = inst[15:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_606 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_48 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [30:0] _next_pc_T_24 = _GEN_31[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 183:40]
  wire [31:0] _next_pc_T_25 = {_GEN_31[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 183:27]
  wire [32:0] _next_reg_1_T_2 = io_now_pc + 32'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 184:31]
  wire [31:0] _next_reg_1_T_3 = io_now_pc + 32'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 184:31]
  wire [3:0] _GEN_2842 = _T_602 ? inst[15:12] : _GEN_2834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2845 = _T_602 ? inst[1:0] : _GEN_2837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2847 = _T_602 | _GEN_2839; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 181:25]
  wire [31:0] _GEN_2848 = _T_602 ? _next_pc_T_23 : _GEN_2840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 183:21]
  wire [31:0] _GEN_2849 = _T_602 ? _next_reg_1_T_1 : _GEN_2832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 184:21]
  wire [2:0] _funct3_T_43 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _ph3_T_2 = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_612 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_1 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_613 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_614 = {2'h1,rs1P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_2850 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_2851 = 5'h1 == _next_reg_T_86 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2852 = 5'h2 == _next_reg_T_86 ? io_now_reg_2 : _GEN_2636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2853 = 5'h3 == _next_reg_T_86 ? io_now_reg_3 : _GEN_2637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2854 = 5'h4 == _next_reg_T_86 ? io_now_reg_4 : _GEN_2638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2855 = 5'h5 == _next_reg_T_86 ? io_now_reg_5 : _GEN_2639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2856 = 5'h6 == _next_reg_T_86 ? io_now_reg_6 : _GEN_2640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2857 = 5'h7 == _next_reg_T_86 ? io_now_reg_7 : _GEN_2641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2858 = 5'h8 == _next_reg_T_86 ? io_now_reg_8 : _GEN_2642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2859 = 5'h9 == _next_reg_T_86 ? io_now_reg_9 : _GEN_2643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2860 = 5'ha == _next_reg_T_86 ? io_now_reg_10 : _GEN_2644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2861 = 5'hb == _next_reg_T_86 ? io_now_reg_11 : _GEN_2645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2862 = 5'hc == _next_reg_T_86 ? io_now_reg_12 : _GEN_2646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2863 = 5'hd == _next_reg_T_86 ? io_now_reg_13 : _GEN_2647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2864 = 5'he == _next_reg_T_86 ? io_now_reg_14 : _GEN_2648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2865 = 5'hf == _next_reg_T_86 ? io_now_reg_15 : _GEN_2649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2866 = 5'h10 == _next_reg_T_86 ? io_now_reg_16 : _GEN_2650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2867 = 5'h11 == _next_reg_T_86 ? io_now_reg_17 : _GEN_2651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2868 = 5'h12 == _next_reg_T_86 ? io_now_reg_18 : _GEN_2652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2869 = 5'h13 == _next_reg_T_86 ? io_now_reg_19 : _GEN_2653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2870 = 5'h14 == _next_reg_T_86 ? io_now_reg_20 : _GEN_2654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2871 = 5'h15 == _next_reg_T_86 ? io_now_reg_21 : _GEN_2655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2872 = 5'h16 == _next_reg_T_86 ? io_now_reg_22 : _GEN_2656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2873 = 5'h17 == _next_reg_T_86 ? io_now_reg_23 : _GEN_2657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2874 = 5'h18 == _next_reg_T_86 ? io_now_reg_24 : _GEN_2658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2875 = 5'h19 == _next_reg_T_86 ? io_now_reg_25 : _GEN_2659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2876 = 5'h1a == _next_reg_T_86 ? io_now_reg_26 : _GEN_2660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2877 = 5'h1b == _next_reg_T_86 ? io_now_reg_27 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2878 = 5'h1c == _next_reg_T_86 ? io_now_reg_28 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2879 = 5'h1d == _next_reg_T_86 ? io_now_reg_29 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2880 = 5'h1e == _next_reg_T_86 ? io_now_reg_30 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _GEN_2881 = 5'h1f == _next_reg_T_86 ? io_now_reg_31 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire [31:0] _now_reg_T_614 = _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:{33,33}]
  wire  _T_615 = _GEN_2666 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:33]
  wire [32:0] _next_pc_T_26 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 191:37]
  wire [31:0] _next_pc_T_27 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 191:37]
  wire  _GEN_2882 = _GEN_2666 == 32'h0 | _GEN_2847; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:42 190:27]
  wire [31:0] _GEN_2883 = _GEN_2666 == 32'h0 ? _T_334 : _GEN_2848; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:42 191:27]
  wire [2:0] _GEN_2885 = _T_608 ? inst[15:13] : _GEN_2826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2886 = _T_608 ? inst[12:10] : _GEN_2808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2888 = _T_608 ? inst[6:2] : _GEN_2586; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2889 = _T_608 ? inst[1:0] : _GEN_2845; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2892 = _T_608 ? _GEN_2882 : _GEN_2847; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24]
  wire [31:0] _GEN_2893 = _T_608 ? _GEN_2883 : _GEN_2848; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24]
  wire [2:0] _funct3_T_44 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _ph3_T_3 = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_621 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_2 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_622 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_623 = {2'h1,rs1P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_2894 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_2895 = 5'h1 == _next_reg_T_86 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2896 = 5'h2 == _next_reg_T_86 ? io_now_reg_2 : _GEN_2636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2897 = 5'h3 == _next_reg_T_86 ? io_now_reg_3 : _GEN_2637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2898 = 5'h4 == _next_reg_T_86 ? io_now_reg_4 : _GEN_2638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2899 = 5'h5 == _next_reg_T_86 ? io_now_reg_5 : _GEN_2639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2900 = 5'h6 == _next_reg_T_86 ? io_now_reg_6 : _GEN_2640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2901 = 5'h7 == _next_reg_T_86 ? io_now_reg_7 : _GEN_2641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2902 = 5'h8 == _next_reg_T_86 ? io_now_reg_8 : _GEN_2642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2903 = 5'h9 == _next_reg_T_86 ? io_now_reg_9 : _GEN_2643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2904 = 5'ha == _next_reg_T_86 ? io_now_reg_10 : _GEN_2644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2905 = 5'hb == _next_reg_T_86 ? io_now_reg_11 : _GEN_2645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2906 = 5'hc == _next_reg_T_86 ? io_now_reg_12 : _GEN_2646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2907 = 5'hd == _next_reg_T_86 ? io_now_reg_13 : _GEN_2647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2908 = 5'he == _next_reg_T_86 ? io_now_reg_14 : _GEN_2648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2909 = 5'hf == _next_reg_T_86 ? io_now_reg_15 : _GEN_2649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2910 = 5'h10 == _next_reg_T_86 ? io_now_reg_16 : _GEN_2650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2911 = 5'h11 == _next_reg_T_86 ? io_now_reg_17 : _GEN_2651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2912 = 5'h12 == _next_reg_T_86 ? io_now_reg_18 : _GEN_2652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2913 = 5'h13 == _next_reg_T_86 ? io_now_reg_19 : _GEN_2653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2914 = 5'h14 == _next_reg_T_86 ? io_now_reg_20 : _GEN_2654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2915 = 5'h15 == _next_reg_T_86 ? io_now_reg_21 : _GEN_2655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2916 = 5'h16 == _next_reg_T_86 ? io_now_reg_22 : _GEN_2656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2917 = 5'h17 == _next_reg_T_86 ? io_now_reg_23 : _GEN_2657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2918 = 5'h18 == _next_reg_T_86 ? io_now_reg_24 : _GEN_2658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2919 = 5'h19 == _next_reg_T_86 ? io_now_reg_25 : _GEN_2659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2920 = 5'h1a == _next_reg_T_86 ? io_now_reg_26 : _GEN_2660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2921 = 5'h1b == _next_reg_T_86 ? io_now_reg_27 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2922 = 5'h1c == _next_reg_T_86 ? io_now_reg_28 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2923 = 5'h1d == _next_reg_T_86 ? io_now_reg_29 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2924 = 5'h1e == _next_reg_T_86 ? io_now_reg_30 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _GEN_2925 = 5'h1f == _next_reg_T_86 ? io_now_reg_31 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire [31:0] _now_reg_T_623 = _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:{33,33}]
  wire  _T_624 = _GEN_2666 != 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:33]
  wire [32:0] _next_pc_T_28 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 199:37]
  wire [31:0] _next_pc_T_29 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 199:37]
  wire  _GEN_2926 = _GEN_2666 != 32'h0 | _GEN_2892; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:42 198:27]
  wire [31:0] _GEN_2927 = _GEN_2666 != 32'h0 ? _T_334 : _GEN_2893; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:42 199:27]
  wire [2:0] _GEN_2929 = _T_617 ? inst[15:13] : _GEN_2885; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2930 = _T_617 ? inst[12:10] : _GEN_2886; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2932 = _T_617 ? inst[6:2] : _GEN_2888; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2933 = _T_617 ? inst[1:0] : _GEN_2889; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2936 = _T_617 ? _GEN_2926 : _GEN_2892; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24]
  wire [31:0] _GEN_2937 = _T_617 ? _GEN_2927 : _GEN_2893; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24]
  wire [2:0] _funct3_T_45 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T_1 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_633 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_3 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_634 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _next_reg_rd_28 = imm; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [31:0] _GEN_2938 = 5'h0 == rd ? imm : _GEN_2710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2939 = 5'h1 == rd ? imm : _GEN_2849; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2940 = 5'h2 == rd ? imm : _GEN_2712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2941 = 5'h3 == rd ? imm : _GEN_2713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2942 = 5'h4 == rd ? imm : _GEN_2714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2943 = 5'h5 == rd ? imm : _GEN_2715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2944 = 5'h6 == rd ? imm : _GEN_2716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2945 = 5'h7 == rd ? imm : _GEN_2717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2946 = 5'h8 == rd ? imm : _GEN_2718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2947 = 5'h9 == rd ? imm : _GEN_2719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2948 = 5'ha == rd ? imm : _GEN_2720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2949 = 5'hb == rd ? imm : _GEN_2721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2950 = 5'hc == rd ? imm : _GEN_2722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2951 = 5'hd == rd ? imm : _GEN_2723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2952 = 5'he == rd ? imm : _GEN_2724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2953 = 5'hf == rd ? imm : _GEN_2725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2954 = 5'h10 == rd ? imm : _GEN_2726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2955 = 5'h11 == rd ? imm : _GEN_2727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2956 = 5'h12 == rd ? imm : _GEN_2728; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2957 = 5'h13 == rd ? imm : _GEN_2729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2958 = 5'h14 == rd ? imm : _GEN_2730; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2959 = 5'h15 == rd ? imm : _GEN_2731; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2960 = 5'h16 == rd ? imm : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2961 = 5'h17 == rd ? imm : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2962 = 5'h18 == rd ? imm : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2963 = 5'h19 == rd ? imm : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2964 = 5'h1a == rd ? imm : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2965 = 5'h1b == rd ? imm : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2966 = 5'h1c == rd ? imm : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2967 = 5'h1d == rd ? imm : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2968 = 5'h1e == rd ? imm : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [31:0] _GEN_2969 = 5'h1f == rd ? imm : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [2:0] _GEN_2971 = _T_629 ? inst[15:13] : _GEN_2929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_2972 = _T_629 ? inst[12] : _GEN_2584; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2974 = _T_629 ? inst[6:2] : _GEN_2932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_2975 = _T_629 ? inst[1:0] : _GEN_2933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2978 = _T_629 ? _GEN_2938 : _GEN_2710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2979 = _T_629 ? _GEN_2939 : _GEN_2849; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2980 = _T_629 ? _GEN_2940 : _GEN_2712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2981 = _T_629 ? _GEN_2941 : _GEN_2713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2982 = _T_629 ? _GEN_2942 : _GEN_2714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2983 = _T_629 ? _GEN_2943 : _GEN_2715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2984 = _T_629 ? _GEN_2944 : _GEN_2716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2985 = _T_629 ? _GEN_2945 : _GEN_2717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2986 = _T_629 ? _GEN_2946 : _GEN_2718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2987 = _T_629 ? _GEN_2947 : _GEN_2719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2988 = _T_629 ? _GEN_2948 : _GEN_2720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2989 = _T_629 ? _GEN_2949 : _GEN_2721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2990 = _T_629 ? _GEN_2950 : _GEN_2722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2991 = _T_629 ? _GEN_2951 : _GEN_2723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2992 = _T_629 ? _GEN_2952 : _GEN_2724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2993 = _T_629 ? _GEN_2953 : _GEN_2725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2994 = _T_629 ? _GEN_2954 : _GEN_2726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2995 = _T_629 ? _GEN_2955 : _GEN_2727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2996 = _T_629 ? _GEN_2956 : _GEN_2728; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2997 = _T_629 ? _GEN_2957 : _GEN_2729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2998 = _T_629 ? _GEN_2958 : _GEN_2730; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_2999 = _T_629 ? _GEN_2959 : _GEN_2731; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3000 = _T_629 ? _GEN_2960 : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3001 = _T_629 ? _GEN_2961 : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3002 = _T_629 ? _GEN_2962 : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3003 = _T_629 ? _GEN_2963 : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3004 = _T_629 ? _GEN_2964 : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3005 = _T_629 ? _GEN_2965 : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3006 = _T_629 ? _GEN_2966 : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3007 = _T_629 ? _GEN_2967 : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3008 = _T_629 ? _GEN_2968 : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [31:0] _GEN_3009 = _T_629 ? _GEN_2969 : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [2:0] _funct3_T_46 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T_2 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_651 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_4 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_652 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _nzimm_C_LUI_T = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_LUI_T_1 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_LUI_T_2 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_LUI_T_3 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_LUI_T_4 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_LUI_T_5 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] nzimm_C_LUI_lo_hi = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [2:0] nzimm_C_LUI_lo = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [1:0] nzimm_C_LUI_hi_hi = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [2:0] nzimm_C_LUI_hi = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [5:0] _nzimm_C_LUI_T_6 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [17:0] _nzimm_C_LUI_T_7 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2],12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  nzimm_C_LUI_signBit = _nzimm_C_LUI_T_7[17]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _nzimm_C_LUI_T_8 = nzimm_C_LUI_signBit; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [13:0] _nzimm_C_LUI_T_9 = nzimm_C_LUI_signBit ? 14'h3fff : 14'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] nzimm_C_LUI = {_nzimm_C_LUI_T_9,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2],12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _next_reg_rd_29 = nzimm_C_LUI; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_3010 = 5'h0 == rd ? nzimm_C_LUI : _GEN_2978; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3011 = 5'h1 == rd ? nzimm_C_LUI : _GEN_2979; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3012 = 5'h2 == rd ? nzimm_C_LUI : _GEN_2980; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3013 = 5'h3 == rd ? nzimm_C_LUI : _GEN_2981; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3014 = 5'h4 == rd ? nzimm_C_LUI : _GEN_2982; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3015 = 5'h5 == rd ? nzimm_C_LUI : _GEN_2983; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3016 = 5'h6 == rd ? nzimm_C_LUI : _GEN_2984; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3017 = 5'h7 == rd ? nzimm_C_LUI : _GEN_2985; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3018 = 5'h8 == rd ? nzimm_C_LUI : _GEN_2986; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3019 = 5'h9 == rd ? nzimm_C_LUI : _GEN_2987; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3020 = 5'ha == rd ? nzimm_C_LUI : _GEN_2988; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3021 = 5'hb == rd ? nzimm_C_LUI : _GEN_2989; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3022 = 5'hc == rd ? nzimm_C_LUI : _GEN_2990; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3023 = 5'hd == rd ? nzimm_C_LUI : _GEN_2991; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3024 = 5'he == rd ? nzimm_C_LUI : _GEN_2992; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3025 = 5'hf == rd ? nzimm_C_LUI : _GEN_2993; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3026 = 5'h10 == rd ? nzimm_C_LUI : _GEN_2994; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3027 = 5'h11 == rd ? nzimm_C_LUI : _GEN_2995; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3028 = 5'h12 == rd ? nzimm_C_LUI : _GEN_2996; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3029 = 5'h13 == rd ? nzimm_C_LUI : _GEN_2997; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3030 = 5'h14 == rd ? nzimm_C_LUI : _GEN_2998; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3031 = 5'h15 == rd ? nzimm_C_LUI : _GEN_2999; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3032 = 5'h16 == rd ? nzimm_C_LUI : _GEN_3000; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3033 = 5'h17 == rd ? nzimm_C_LUI : _GEN_3001; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3034 = 5'h18 == rd ? nzimm_C_LUI : _GEN_3002; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3035 = 5'h19 == rd ? nzimm_C_LUI : _GEN_3003; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3036 = 5'h1a == rd ? nzimm_C_LUI : _GEN_3004; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3037 = 5'h1b == rd ? nzimm_C_LUI : _GEN_3005; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3038 = 5'h1c == rd ? nzimm_C_LUI : _GEN_3006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3039 = 5'h1d == rd ? nzimm_C_LUI : _GEN_3007; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3040 = 5'h1e == rd ? nzimm_C_LUI : _GEN_3008; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [31:0] _GEN_3041 = 5'h1f == rd ? nzimm_C_LUI : _GEN_3009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [2:0] _GEN_3043 = _T_647 ? inst[15:13] : _GEN_2971; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_3044 = _T_647 ? inst[12] : _GEN_2972; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3046 = _T_647 ? inst[6:2] : _GEN_2974; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3047 = _T_647 ? inst[1:0] : _GEN_2975; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3049 = _T_647 ? _GEN_3010 : _GEN_2978; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3050 = _T_647 ? _GEN_3011 : _GEN_2979; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3051 = _T_647 ? _GEN_3012 : _GEN_2980; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3052 = _T_647 ? _GEN_3013 : _GEN_2981; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3053 = _T_647 ? _GEN_3014 : _GEN_2982; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3054 = _T_647 ? _GEN_3015 : _GEN_2983; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3055 = _T_647 ? _GEN_3016 : _GEN_2984; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3056 = _T_647 ? _GEN_3017 : _GEN_2985; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3057 = _T_647 ? _GEN_3018 : _GEN_2986; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3058 = _T_647 ? _GEN_3019 : _GEN_2987; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3059 = _T_647 ? _GEN_3020 : _GEN_2988; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3060 = _T_647 ? _GEN_3021 : _GEN_2989; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3061 = _T_647 ? _GEN_3022 : _GEN_2990; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3062 = _T_647 ? _GEN_3023 : _GEN_2991; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3063 = _T_647 ? _GEN_3024 : _GEN_2992; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3064 = _T_647 ? _GEN_3025 : _GEN_2993; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3065 = _T_647 ? _GEN_3026 : _GEN_2994; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3066 = _T_647 ? _GEN_3027 : _GEN_2995; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3067 = _T_647 ? _GEN_3028 : _GEN_2996; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3068 = _T_647 ? _GEN_3029 : _GEN_2997; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3069 = _T_647 ? _GEN_3030 : _GEN_2998; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3070 = _T_647 ? _GEN_3031 : _GEN_2999; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3071 = _T_647 ? _GEN_3032 : _GEN_3000; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3072 = _T_647 ? _GEN_3033 : _GEN_3001; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3073 = _T_647 ? _GEN_3034 : _GEN_3002; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3074 = _T_647 ? _GEN_3035 : _GEN_3003; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3075 = _T_647 ? _GEN_3036 : _GEN_3004; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3076 = _T_647 ? _GEN_3037 : _GEN_3005; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3077 = _T_647 ? _GEN_3038 : _GEN_3006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3078 = _T_647 ? _GEN_3039 : _GEN_3007; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3079 = _T_647 ? _GEN_3040 : _GEN_3008; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [31:0] _GEN_3080 = _T_647 ? _GEN_3041 : _GEN_3009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [2:0] _funct3_T_47 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T_3 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_666 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_5 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_667 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _nzimm_C_ADDI_T = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _nzimm_C_ADDI_T_1 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _nzimm_C_ADDI_T_2 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _nzimm_C_ADDI_T_3 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _nzimm_C_ADDI_T_4 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire  _nzimm_C_ADDI_T_5 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:32]
  wire [1:0] nzimm_C_ADDI_lo_hi = {inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [2:0] nzimm_C_ADDI_lo = {inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [1:0] nzimm_C_ADDI_hi_hi = {inst[12],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [2:0] nzimm_C_ADDI_hi = {inst[12],inst[6],inst[5]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire [5:0] _nzimm_C_ADDI_T_6 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  nzimm_C_ADDI_signBit = _imm_T_227[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _nzimm_C_ADDI_T_7 = imm_signBit_35; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [25:0] _nzimm_C_ADDI_T_8 = imm_signBit_35 ? 26'h3ffffff : 26'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] nzimm_C_ADDI = {_imm_T_229,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_3081 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3082 = 5'h1 == rd ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3083 = 5'h2 == rd ? io_now_reg_2 : _GEN_3082; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3084 = 5'h3 == rd ? io_now_reg_3 : _GEN_3083; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3085 = 5'h4 == rd ? io_now_reg_4 : _GEN_3084; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3086 = 5'h5 == rd ? io_now_reg_5 : _GEN_3085; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3087 = 5'h6 == rd ? io_now_reg_6 : _GEN_3086; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3088 = 5'h7 == rd ? io_now_reg_7 : _GEN_3087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3089 = 5'h8 == rd ? io_now_reg_8 : _GEN_3088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3090 = 5'h9 == rd ? io_now_reg_9 : _GEN_3089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3091 = 5'ha == rd ? io_now_reg_10 : _GEN_3090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3092 = 5'hb == rd ? io_now_reg_11 : _GEN_3091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3093 = 5'hc == rd ? io_now_reg_12 : _GEN_3092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3094 = 5'hd == rd ? io_now_reg_13 : _GEN_3093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3095 = 5'he == rd ? io_now_reg_14 : _GEN_3094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3096 = 5'hf == rd ? io_now_reg_15 : _GEN_3095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3097 = 5'h10 == rd ? io_now_reg_16 : _GEN_3096; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3098 = 5'h11 == rd ? io_now_reg_17 : _GEN_3097; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3099 = 5'h12 == rd ? io_now_reg_18 : _GEN_3098; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3100 = 5'h13 == rd ? io_now_reg_19 : _GEN_3099; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3101 = 5'h14 == rd ? io_now_reg_20 : _GEN_3100; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3102 = 5'h15 == rd ? io_now_reg_21 : _GEN_3101; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3103 = 5'h16 == rd ? io_now_reg_22 : _GEN_3102; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3104 = 5'h17 == rd ? io_now_reg_23 : _GEN_3103; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3105 = 5'h18 == rd ? io_now_reg_24 : _GEN_3104; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3106 = 5'h19 == rd ? io_now_reg_25 : _GEN_3105; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3107 = 5'h1a == rd ? io_now_reg_26 : _GEN_3106; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3108 = 5'h1b == rd ? io_now_reg_27 : _GEN_3107; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3109 = 5'h1c == rd ? io_now_reg_28 : _GEN_3108; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3110 = 5'h1d == rd ? io_now_reg_29 : _GEN_3109; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3111 = 5'h1e == rd ? io_now_reg_30 : _GEN_3110; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _GEN_3112 = 5'h1f == rd ? io_now_reg_31 : _GEN_3111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _now_reg_rd = 5'h1f == rd ? io_now_reg_31 : _GEN_3111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [32:0] _next_reg_T_93 = _GEN_3112 + _imm_T_230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:35]
  wire [31:0] _next_reg_T_94 = _GEN_3112 + _imm_T_230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:35]
  wire [31:0] _next_reg_rd_30 = _GEN_3112 + _imm_T_230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:35]
  wire [31:0] _GEN_3113 = 5'h0 == rd ? _next_reg_T_94 : _GEN_3049; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3114 = 5'h1 == rd ? _next_reg_T_94 : _GEN_3050; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3115 = 5'h2 == rd ? _next_reg_T_94 : _GEN_3051; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3116 = 5'h3 == rd ? _next_reg_T_94 : _GEN_3052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3117 = 5'h4 == rd ? _next_reg_T_94 : _GEN_3053; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3118 = 5'h5 == rd ? _next_reg_T_94 : _GEN_3054; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3119 = 5'h6 == rd ? _next_reg_T_94 : _GEN_3055; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3120 = 5'h7 == rd ? _next_reg_T_94 : _GEN_3056; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3121 = 5'h8 == rd ? _next_reg_T_94 : _GEN_3057; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3122 = 5'h9 == rd ? _next_reg_T_94 : _GEN_3058; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3123 = 5'ha == rd ? _next_reg_T_94 : _GEN_3059; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3124 = 5'hb == rd ? _next_reg_T_94 : _GEN_3060; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3125 = 5'hc == rd ? _next_reg_T_94 : _GEN_3061; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3126 = 5'hd == rd ? _next_reg_T_94 : _GEN_3062; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3127 = 5'he == rd ? _next_reg_T_94 : _GEN_3063; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3128 = 5'hf == rd ? _next_reg_T_94 : _GEN_3064; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3129 = 5'h10 == rd ? _next_reg_T_94 : _GEN_3065; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3130 = 5'h11 == rd ? _next_reg_T_94 : _GEN_3066; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3131 = 5'h12 == rd ? _next_reg_T_94 : _GEN_3067; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3132 = 5'h13 == rd ? _next_reg_T_94 : _GEN_3068; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3133 = 5'h14 == rd ? _next_reg_T_94 : _GEN_3069; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3134 = 5'h15 == rd ? _next_reg_T_94 : _GEN_3070; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3135 = 5'h16 == rd ? _next_reg_T_94 : _GEN_3071; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3136 = 5'h17 == rd ? _next_reg_T_94 : _GEN_3072; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3137 = 5'h18 == rd ? _next_reg_T_94 : _GEN_3073; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3138 = 5'h19 == rd ? _next_reg_T_94 : _GEN_3074; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3139 = 5'h1a == rd ? _next_reg_T_94 : _GEN_3075; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3140 = 5'h1b == rd ? _next_reg_T_94 : _GEN_3076; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3141 = 5'h1c == rd ? _next_reg_T_94 : _GEN_3077; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3142 = 5'h1d == rd ? _next_reg_T_94 : _GEN_3078; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3143 = 5'h1e == rd ? _next_reg_T_94 : _GEN_3079; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [31:0] _GEN_3144 = 5'h1f == rd ? _next_reg_T_94 : _GEN_3080; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [2:0] _GEN_3146 = _T_662 ? inst[15:13] : _GEN_3043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_3147 = _T_662 ? inst[12] : _GEN_3044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3149 = _T_662 ? inst[6:2] : _GEN_3046; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3150 = _T_662 ? inst[1:0] : _GEN_3047; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3152 = _T_662 ? _GEN_3113 : _GEN_3049; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3153 = _T_662 ? _GEN_3114 : _GEN_3050; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3154 = _T_662 ? _GEN_3115 : _GEN_3051; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3155 = _T_662 ? _GEN_3116 : _GEN_3052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3156 = _T_662 ? _GEN_3117 : _GEN_3053; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3157 = _T_662 ? _GEN_3118 : _GEN_3054; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3158 = _T_662 ? _GEN_3119 : _GEN_3055; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3159 = _T_662 ? _GEN_3120 : _GEN_3056; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3160 = _T_662 ? _GEN_3121 : _GEN_3057; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3161 = _T_662 ? _GEN_3122 : _GEN_3058; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3162 = _T_662 ? _GEN_3123 : _GEN_3059; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3163 = _T_662 ? _GEN_3124 : _GEN_3060; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3164 = _T_662 ? _GEN_3125 : _GEN_3061; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3165 = _T_662 ? _GEN_3126 : _GEN_3062; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3166 = _T_662 ? _GEN_3127 : _GEN_3063; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3167 = _T_662 ? _GEN_3128 : _GEN_3064; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3168 = _T_662 ? _GEN_3129 : _GEN_3065; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3169 = _T_662 ? _GEN_3130 : _GEN_3066; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3170 = _T_662 ? _GEN_3131 : _GEN_3067; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3171 = _T_662 ? _GEN_3132 : _GEN_3068; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3172 = _T_662 ? _GEN_3133 : _GEN_3069; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3173 = _T_662 ? _GEN_3134 : _GEN_3070; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3174 = _T_662 ? _GEN_3135 : _GEN_3071; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3175 = _T_662 ? _GEN_3136 : _GEN_3072; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3176 = _T_662 ? _GEN_3137 : _GEN_3073; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3177 = _T_662 ? _GEN_3138 : _GEN_3074; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3178 = _T_662 ? _GEN_3139 : _GEN_3075; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3179 = _T_662 ? _GEN_3140 : _GEN_3076; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3180 = _T_662 ? _GEN_3141 : _GEN_3077; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3181 = _T_662 ? _GEN_3142 : _GEN_3078; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3182 = _T_662 ? _GEN_3143 : _GEN_3079; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [31:0] _GEN_3183 = _T_662 ? _GEN_3144 : _GEN_3080; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [2:0] _funct3_T_48 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T_4 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_678 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_6 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_679 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _nzimm_C_ADDI16SP_T = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI16SP_T_1 = inst[4]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI16SP_T_2 = inst[3]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI16SP_T_3 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI16SP_T_4 = inst[2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI16SP_T_5 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] nzimm_C_ADDI16SP_lo_hi = {inst[5],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [2:0] nzimm_C_ADDI16SP_lo = {inst[5],inst[2],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [1:0] nzimm_C_ADDI16SP_hi_hi = {inst[12],inst[4]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [2:0] nzimm_C_ADDI16SP_hi = {inst[12],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [5:0] _nzimm_C_ADDI16SP_T_6 = {inst[12],inst[4],inst[3],inst[5],inst[2],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [9:0] _nzimm_C_ADDI16SP_T_7 = {inst[12],inst[4],inst[3],inst[5],inst[2],inst[6],4'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  nzimm_C_ADDI16SP_signBit = _nzimm_C_ADDI16SP_T_7[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _nzimm_C_ADDI16SP_T_8 = nzimm_C_ADDI16SP_signBit; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [21:0] _nzimm_C_ADDI16SP_T_9 = nzimm_C_ADDI16SP_signBit ? 22'h3fffff : 22'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] nzimm_C_ADDI16SP = {_nzimm_C_ADDI16SP_T_9,inst[12],inst[4],inst[3],inst[5],inst[2],inst[6],4'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [32:0] _next_reg_2_T = io_now_reg_2 + nzimm_C_ADDI16SP; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 223:37]
  wire [31:0] _next_reg_2_T_1 = io_now_reg_2 + nzimm_C_ADDI16SP; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 223:37]
  wire [2:0] _GEN_3185 = _T_674 ? inst[15:13] : _GEN_3146; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_3186 = _T_674 ? inst[12] : _GEN_3147; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3188 = _T_674 ? inst[6:2] : _GEN_3149; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3189 = _T_674 ? inst[1:0] : _GEN_3150; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3191 = _T_674 ? _next_reg_2_T_1 : _GEN_3154; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 223:21]
  wire [2:0] _funct3_T_49 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [7:0] _ph8_T = inst[12:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_688 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _nzimm_C_ADDI4SPN_T = inst[10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_1 = inst[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_2 = inst[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_3 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_4 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_5 = inst[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_6 = inst[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire  _nzimm_C_ADDI4SPN_T_7 = inst[6]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:36]
  wire [1:0] nzimm_C_ADDI4SPN_lo_lo = {inst[5],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [1:0] nzimm_C_ADDI4SPN_lo_hi = {inst[12],inst[11]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [3:0] nzimm_C_ADDI4SPN_lo = {inst[12],inst[11],inst[5],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [1:0] nzimm_C_ADDI4SPN_hi_lo = {inst[8],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [1:0] nzimm_C_ADDI4SPN_hi_hi = {inst[10],inst[9]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [3:0] nzimm_C_ADDI4SPN_hi = {inst[10],inst[9],inst[8],inst[7]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [7:0] _nzimm_C_ADDI4SPN_T_8 = {inst[10],inst[9],inst[8],inst[7],inst[12],inst[11],inst[5],inst[6]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [9:0] _nzimm_C_ADDI4SPN_T_9 = {inst[10],inst[9],inst[8],inst[7],inst[12],inst[11],inst[5],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire [31:0] nzimm_C_ADDI4SPN = {22'h0,inst[10],inst[9],inst[8],inst[7],inst[12],inst[11],inst[5],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [4:0] _T_689 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [32:0] _next_reg_T_95 = io_now_reg_2 + nzimm_C_ADDI4SPN; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:44]
  wire [31:0] _next_reg_T_96 = io_now_reg_2 + nzimm_C_ADDI4SPN; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:44]
  wire [31:0] _next_reg_T_689 = io_now_reg_2 + nzimm_C_ADDI4SPN; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:44]
  wire [31:0] _GEN_3192 = 5'h0 == _T_565 ? _next_reg_T_96 : _GEN_3152; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3193 = 5'h1 == _T_565 ? _next_reg_T_96 : _GEN_3153; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3194 = 5'h2 == _T_565 ? _next_reg_T_96 : _GEN_3191; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3195 = 5'h3 == _T_565 ? _next_reg_T_96 : _GEN_3155; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3196 = 5'h4 == _T_565 ? _next_reg_T_96 : _GEN_3156; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3197 = 5'h5 == _T_565 ? _next_reg_T_96 : _GEN_3157; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3198 = 5'h6 == _T_565 ? _next_reg_T_96 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3199 = 5'h7 == _T_565 ? _next_reg_T_96 : _GEN_3159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3200 = 5'h8 == _T_565 ? _next_reg_T_96 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3201 = 5'h9 == _T_565 ? _next_reg_T_96 : _GEN_3161; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3202 = 5'ha == _T_565 ? _next_reg_T_96 : _GEN_3162; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3203 = 5'hb == _T_565 ? _next_reg_T_96 : _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3204 = 5'hc == _T_565 ? _next_reg_T_96 : _GEN_3164; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3205 = 5'hd == _T_565 ? _next_reg_T_96 : _GEN_3165; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3206 = 5'he == _T_565 ? _next_reg_T_96 : _GEN_3166; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3207 = 5'hf == _T_565 ? _next_reg_T_96 : _GEN_3167; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3208 = 5'h10 == _T_565 ? _next_reg_T_96 : _GEN_3168; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3209 = 5'h11 == _T_565 ? _next_reg_T_96 : _GEN_3169; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3210 = 5'h12 == _T_565 ? _next_reg_T_96 : _GEN_3170; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3211 = 5'h13 == _T_565 ? _next_reg_T_96 : _GEN_3171; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3212 = 5'h14 == _T_565 ? _next_reg_T_96 : _GEN_3172; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3213 = 5'h15 == _T_565 ? _next_reg_T_96 : _GEN_3173; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3214 = 5'h16 == _T_565 ? _next_reg_T_96 : _GEN_3174; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3215 = 5'h17 == _T_565 ? _next_reg_T_96 : _GEN_3175; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3216 = 5'h18 == _T_565 ? _next_reg_T_96 : _GEN_3176; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3217 = 5'h19 == _T_565 ? _next_reg_T_96 : _GEN_3177; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3218 = 5'h1a == _T_565 ? _next_reg_T_96 : _GEN_3178; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3219 = 5'h1b == _T_565 ? _next_reg_T_96 : _GEN_3179; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3220 = 5'h1c == _T_565 ? _next_reg_T_96 : _GEN_3180; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3221 = 5'h1d == _T_565 ? _next_reg_T_96 : _GEN_3181; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3222 = 5'h1e == _T_565 ? _next_reg_T_96 : _GEN_3182; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [31:0] _GEN_3223 = 5'h1f == _T_565 ? _next_reg_T_96 : _GEN_3183; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [2:0] _GEN_3225 = _T_684 ? inst[15:13] : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [7:0] _GEN_3226 = _T_684 ? inst[12:5] : 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 105:22]
  wire [1:0] _GEN_3228 = _T_684 ? inst[1:0] : _GEN_3189; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3229 = _T_684 ? _GEN_3192 : _GEN_3152; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3230 = _T_684 ? _GEN_3193 : _GEN_3153; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3231 = _T_684 ? _GEN_3194 : _GEN_3191; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3232 = _T_684 ? _GEN_3195 : _GEN_3155; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3233 = _T_684 ? _GEN_3196 : _GEN_3156; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3234 = _T_684 ? _GEN_3197 : _GEN_3157; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3235 = _T_684 ? _GEN_3198 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3236 = _T_684 ? _GEN_3199 : _GEN_3159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3237 = _T_684 ? _GEN_3200 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3238 = _T_684 ? _GEN_3201 : _GEN_3161; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3239 = _T_684 ? _GEN_3202 : _GEN_3162; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3240 = _T_684 ? _GEN_3203 : _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3241 = _T_684 ? _GEN_3204 : _GEN_3164; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3242 = _T_684 ? _GEN_3205 : _GEN_3165; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3243 = _T_684 ? _GEN_3206 : _GEN_3166; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3244 = _T_684 ? _GEN_3207 : _GEN_3167; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3245 = _T_684 ? _GEN_3208 : _GEN_3168; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3246 = _T_684 ? _GEN_3209 : _GEN_3169; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3247 = _T_684 ? _GEN_3210 : _GEN_3170; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3248 = _T_684 ? _GEN_3211 : _GEN_3171; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3249 = _T_684 ? _GEN_3212 : _GEN_3172; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3250 = _T_684 ? _GEN_3213 : _GEN_3173; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3251 = _T_684 ? _GEN_3214 : _GEN_3174; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3252 = _T_684 ? _GEN_3215 : _GEN_3175; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3253 = _T_684 ? _GEN_3216 : _GEN_3176; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3254 = _T_684 ? _GEN_3217 : _GEN_3177; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3255 = _T_684 ? _GEN_3218 : _GEN_3178; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3256 = _T_684 ? _GEN_3219 : _GEN_3179; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3257 = _T_684 ? _GEN_3220 : _GEN_3180; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3258 = _T_684 ? _GEN_3221 : _GEN_3181; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3259 = _T_684 ? _GEN_3222 : _GEN_3182; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [31:0] _GEN_3260 = _T_684 ? _GEN_3223 : _GEN_3183; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [2:0] _funct3_T_50 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T_5 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_706 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_7 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_707 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [5:0] _next_reg_T_97 = imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:41]
  wire [31:0] _now_reg_rd_0 = 5'h1f == rd ? io_now_reg_31 : _GEN_3111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [94:0] _GEN_6219 = {{63'd0}, _GEN_3112}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:35]
  wire [94:0] _next_reg_T_98 = _GEN_6219 << imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:35]
  wire [31:0] _next_reg_rd_31 = _next_reg_T_98[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3261 = 5'h0 == rd ? _next_reg_T_98[31:0] : _GEN_3229; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3262 = 5'h1 == rd ? _next_reg_T_98[31:0] : _GEN_3230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3263 = 5'h2 == rd ? _next_reg_T_98[31:0] : _GEN_3231; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3264 = 5'h3 == rd ? _next_reg_T_98[31:0] : _GEN_3232; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3265 = 5'h4 == rd ? _next_reg_T_98[31:0] : _GEN_3233; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3266 = 5'h5 == rd ? _next_reg_T_98[31:0] : _GEN_3234; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3267 = 5'h6 == rd ? _next_reg_T_98[31:0] : _GEN_3235; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3268 = 5'h7 == rd ? _next_reg_T_98[31:0] : _GEN_3236; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3269 = 5'h8 == rd ? _next_reg_T_98[31:0] : _GEN_3237; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3270 = 5'h9 == rd ? _next_reg_T_98[31:0] : _GEN_3238; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3271 = 5'ha == rd ? _next_reg_T_98[31:0] : _GEN_3239; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3272 = 5'hb == rd ? _next_reg_T_98[31:0] : _GEN_3240; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3273 = 5'hc == rd ? _next_reg_T_98[31:0] : _GEN_3241; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3274 = 5'hd == rd ? _next_reg_T_98[31:0] : _GEN_3242; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3275 = 5'he == rd ? _next_reg_T_98[31:0] : _GEN_3243; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3276 = 5'hf == rd ? _next_reg_T_98[31:0] : _GEN_3244; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3277 = 5'h10 == rd ? _next_reg_T_98[31:0] : _GEN_3245; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3278 = 5'h11 == rd ? _next_reg_T_98[31:0] : _GEN_3246; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3279 = 5'h12 == rd ? _next_reg_T_98[31:0] : _GEN_3247; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3280 = 5'h13 == rd ? _next_reg_T_98[31:0] : _GEN_3248; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3281 = 5'h14 == rd ? _next_reg_T_98[31:0] : _GEN_3249; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3282 = 5'h15 == rd ? _next_reg_T_98[31:0] : _GEN_3250; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3283 = 5'h16 == rd ? _next_reg_T_98[31:0] : _GEN_3251; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3284 = 5'h17 == rd ? _next_reg_T_98[31:0] : _GEN_3252; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3285 = 5'h18 == rd ? _next_reg_T_98[31:0] : _GEN_3253; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3286 = 5'h19 == rd ? _next_reg_T_98[31:0] : _GEN_3254; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3287 = 5'h1a == rd ? _next_reg_T_98[31:0] : _GEN_3255; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3288 = 5'h1b == rd ? _next_reg_T_98[31:0] : _GEN_3256; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3289 = 5'h1c == rd ? _next_reg_T_98[31:0] : _GEN_3257; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3290 = 5'h1d == rd ? _next_reg_T_98[31:0] : _GEN_3258; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3291 = 5'h1e == rd ? _next_reg_T_98[31:0] : _GEN_3259; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [31:0] _GEN_3292 = 5'h1f == rd ? _next_reg_T_98[31:0] : _GEN_3260; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [2:0] _GEN_3294 = _T_702 ? inst[15:13] : _GEN_3225; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_3295 = _T_702 ? inst[12] : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3297 = _T_702 ? inst[6:2] : _GEN_3188; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3298 = _T_702 ? inst[1:0] : _GEN_3228; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3301 = _T_702 ? _GEN_3261 : _GEN_3229; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3302 = _T_702 ? _GEN_3262 : _GEN_3230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3303 = _T_702 ? _GEN_3263 : _GEN_3231; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3304 = _T_702 ? _GEN_3264 : _GEN_3232; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3305 = _T_702 ? _GEN_3265 : _GEN_3233; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3306 = _T_702 ? _GEN_3266 : _GEN_3234; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3307 = _T_702 ? _GEN_3267 : _GEN_3235; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3308 = _T_702 ? _GEN_3268 : _GEN_3236; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3309 = _T_702 ? _GEN_3269 : _GEN_3237; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3310 = _T_702 ? _GEN_3270 : _GEN_3238; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3311 = _T_702 ? _GEN_3271 : _GEN_3239; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3312 = _T_702 ? _GEN_3272 : _GEN_3240; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3313 = _T_702 ? _GEN_3273 : _GEN_3241; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3314 = _T_702 ? _GEN_3274 : _GEN_3242; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3315 = _T_702 ? _GEN_3275 : _GEN_3243; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3316 = _T_702 ? _GEN_3276 : _GEN_3244; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3317 = _T_702 ? _GEN_3277 : _GEN_3245; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3318 = _T_702 ? _GEN_3278 : _GEN_3246; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3319 = _T_702 ? _GEN_3279 : _GEN_3247; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3320 = _T_702 ? _GEN_3280 : _GEN_3248; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3321 = _T_702 ? _GEN_3281 : _GEN_3249; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3322 = _T_702 ? _GEN_3282 : _GEN_3250; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3323 = _T_702 ? _GEN_3283 : _GEN_3251; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3324 = _T_702 ? _GEN_3284 : _GEN_3252; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3325 = _T_702 ? _GEN_3285 : _GEN_3253; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3326 = _T_702 ? _GEN_3286 : _GEN_3254; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3327 = _T_702 ? _GEN_3287 : _GEN_3255; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3328 = _T_702 ? _GEN_3288 : _GEN_3256; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3329 = _T_702 ? _GEN_3289 : _GEN_3257; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3330 = _T_702 ? _GEN_3290 : _GEN_3258; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3331 = _T_702 ? _GEN_3291 : _GEN_3259; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [31:0] _GEN_3332 = _T_702 ? _GEN_3292 : _GEN_3260; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [2:0] _funct3_T_51 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _ph3_T_4 = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_721 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_8 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_722 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_723 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_99 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [5:0] _next_reg_T_100 = imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:57]
  wire [31:0] _GEN_3333 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3334 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3335 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3336 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3337 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3338 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3339 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3340 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3341 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3342 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3343 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3344 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3345 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3346 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3347 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3348 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3349 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3350 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3351 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3352 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3353 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3354 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3355 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3356 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3357 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3358 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3359 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3360 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3361 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3362 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3363 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _GEN_3364 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _now_reg_next_reg_T_99 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [31:0] _next_reg_T_101 = _GEN_3364 >> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:51]
  wire [31:0] _next_reg_T_723 = _GEN_3364 >> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:51]
  wire [31:0] _GEN_3365 = 5'h0 == _T_565 ? _next_reg_T_101 : _GEN_3301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3366 = 5'h1 == _T_565 ? _next_reg_T_101 : _GEN_3302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3367 = 5'h2 == _T_565 ? _next_reg_T_101 : _GEN_3303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3368 = 5'h3 == _T_565 ? _next_reg_T_101 : _GEN_3304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3369 = 5'h4 == _T_565 ? _next_reg_T_101 : _GEN_3305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3370 = 5'h5 == _T_565 ? _next_reg_T_101 : _GEN_3306; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3371 = 5'h6 == _T_565 ? _next_reg_T_101 : _GEN_3307; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3372 = 5'h7 == _T_565 ? _next_reg_T_101 : _GEN_3308; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3373 = 5'h8 == _T_565 ? _next_reg_T_101 : _GEN_3309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3374 = 5'h9 == _T_565 ? _next_reg_T_101 : _GEN_3310; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3375 = 5'ha == _T_565 ? _next_reg_T_101 : _GEN_3311; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3376 = 5'hb == _T_565 ? _next_reg_T_101 : _GEN_3312; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3377 = 5'hc == _T_565 ? _next_reg_T_101 : _GEN_3313; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3378 = 5'hd == _T_565 ? _next_reg_T_101 : _GEN_3314; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3379 = 5'he == _T_565 ? _next_reg_T_101 : _GEN_3315; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3380 = 5'hf == _T_565 ? _next_reg_T_101 : _GEN_3316; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3381 = 5'h10 == _T_565 ? _next_reg_T_101 : _GEN_3317; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3382 = 5'h11 == _T_565 ? _next_reg_T_101 : _GEN_3318; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3383 = 5'h12 == _T_565 ? _next_reg_T_101 : _GEN_3319; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3384 = 5'h13 == _T_565 ? _next_reg_T_101 : _GEN_3320; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3385 = 5'h14 == _T_565 ? _next_reg_T_101 : _GEN_3321; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3386 = 5'h15 == _T_565 ? _next_reg_T_101 : _GEN_3322; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3387 = 5'h16 == _T_565 ? _next_reg_T_101 : _GEN_3323; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3388 = 5'h17 == _T_565 ? _next_reg_T_101 : _GEN_3324; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3389 = 5'h18 == _T_565 ? _next_reg_T_101 : _GEN_3325; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3390 = 5'h19 == _T_565 ? _next_reg_T_101 : _GEN_3326; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3391 = 5'h1a == _T_565 ? _next_reg_T_101 : _GEN_3327; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3392 = 5'h1b == _T_565 ? _next_reg_T_101 : _GEN_3328; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3393 = 5'h1c == _T_565 ? _next_reg_T_101 : _GEN_3329; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3394 = 5'h1d == _T_565 ? _next_reg_T_101 : _GEN_3330; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3395 = 5'h1e == _T_565 ? _next_reg_T_101 : _GEN_3331; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [31:0] _GEN_3396 = 5'h1f == _T_565 ? _next_reg_T_101 : _GEN_3332; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [2:0] _GEN_3398 = _T_717 ? inst[15:13] : _GEN_3294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3399 = _T_717 ? inst[12:10] : _GEN_2930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3401 = _T_717 ? inst[6:2] : _GEN_3297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3402 = _T_717 ? inst[1:0] : _GEN_3298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3405 = _T_717 ? _GEN_3365 : _GEN_3301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3406 = _T_717 ? _GEN_3366 : _GEN_3302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3407 = _T_717 ? _GEN_3367 : _GEN_3303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3408 = _T_717 ? _GEN_3368 : _GEN_3304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3409 = _T_717 ? _GEN_3369 : _GEN_3305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3410 = _T_717 ? _GEN_3370 : _GEN_3306; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3411 = _T_717 ? _GEN_3371 : _GEN_3307; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3412 = _T_717 ? _GEN_3372 : _GEN_3308; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3413 = _T_717 ? _GEN_3373 : _GEN_3309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3414 = _T_717 ? _GEN_3374 : _GEN_3310; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3415 = _T_717 ? _GEN_3375 : _GEN_3311; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3416 = _T_717 ? _GEN_3376 : _GEN_3312; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3417 = _T_717 ? _GEN_3377 : _GEN_3313; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3418 = _T_717 ? _GEN_3378 : _GEN_3314; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3419 = _T_717 ? _GEN_3379 : _GEN_3315; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3420 = _T_717 ? _GEN_3380 : _GEN_3316; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3421 = _T_717 ? _GEN_3381 : _GEN_3317; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3422 = _T_717 ? _GEN_3382 : _GEN_3318; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3423 = _T_717 ? _GEN_3383 : _GEN_3319; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3424 = _T_717 ? _GEN_3384 : _GEN_3320; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3425 = _T_717 ? _GEN_3385 : _GEN_3321; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3426 = _T_717 ? _GEN_3386 : _GEN_3322; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3427 = _T_717 ? _GEN_3387 : _GEN_3323; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3428 = _T_717 ? _GEN_3388 : _GEN_3324; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3429 = _T_717 ? _GEN_3389 : _GEN_3325; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3430 = _T_717 ? _GEN_3390 : _GEN_3326; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3431 = _T_717 ? _GEN_3391 : _GEN_3327; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3432 = _T_717 ? _GEN_3392 : _GEN_3328; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3433 = _T_717 ? _GEN_3393 : _GEN_3329; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3434 = _T_717 ? _GEN_3394 : _GEN_3330; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3435 = _T_717 ? _GEN_3395 : _GEN_3331; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [31:0] _GEN_3436 = _T_717 ? _GEN_3396 : _GEN_3332; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [2:0] _funct3_T_52 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _ph3_T_5 = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_737 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_9 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_738 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_739 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_102 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_3437 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3438 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3439 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3440 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3441 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3442 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3443 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3444 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3445 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3446 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3447 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3448 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3449 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3450 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3451 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3452 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3453 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3454 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3455 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3456 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3457 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3458 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3459 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3460 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3461 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3462 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3463 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3464 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3465 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3466 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3467 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _GEN_3468 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _now_reg_next_reg_T_102 = _GEN_3364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{52,52}]
  wire [31:0] _next_reg_T_103 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:52]
  wire [5:0] _next_reg_T_104 = imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:65]
  wire [31:0] _next_reg_T_105 = $signed(_next_reg_T_103) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:59]
  wire [31:0] _next_reg_T_106 = $signed(_next_reg_T_103) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:73]
  wire [31:0] _next_reg_T_739 = $signed(_next_reg_T_103) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:73]
  wire [31:0] _GEN_3469 = 5'h0 == _T_565 ? _next_reg_T_106 : _GEN_3405; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3470 = 5'h1 == _T_565 ? _next_reg_T_106 : _GEN_3406; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3471 = 5'h2 == _T_565 ? _next_reg_T_106 : _GEN_3407; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3472 = 5'h3 == _T_565 ? _next_reg_T_106 : _GEN_3408; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3473 = 5'h4 == _T_565 ? _next_reg_T_106 : _GEN_3409; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3474 = 5'h5 == _T_565 ? _next_reg_T_106 : _GEN_3410; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3475 = 5'h6 == _T_565 ? _next_reg_T_106 : _GEN_3411; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3476 = 5'h7 == _T_565 ? _next_reg_T_106 : _GEN_3412; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3477 = 5'h8 == _T_565 ? _next_reg_T_106 : _GEN_3413; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3478 = 5'h9 == _T_565 ? _next_reg_T_106 : _GEN_3414; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3479 = 5'ha == _T_565 ? _next_reg_T_106 : _GEN_3415; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3480 = 5'hb == _T_565 ? _next_reg_T_106 : _GEN_3416; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3481 = 5'hc == _T_565 ? _next_reg_T_106 : _GEN_3417; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3482 = 5'hd == _T_565 ? _next_reg_T_106 : _GEN_3418; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3483 = 5'he == _T_565 ? _next_reg_T_106 : _GEN_3419; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3484 = 5'hf == _T_565 ? _next_reg_T_106 : _GEN_3420; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3485 = 5'h10 == _T_565 ? _next_reg_T_106 : _GEN_3421; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3486 = 5'h11 == _T_565 ? _next_reg_T_106 : _GEN_3422; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3487 = 5'h12 == _T_565 ? _next_reg_T_106 : _GEN_3423; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3488 = 5'h13 == _T_565 ? _next_reg_T_106 : _GEN_3424; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3489 = 5'h14 == _T_565 ? _next_reg_T_106 : _GEN_3425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3490 = 5'h15 == _T_565 ? _next_reg_T_106 : _GEN_3426; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3491 = 5'h16 == _T_565 ? _next_reg_T_106 : _GEN_3427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3492 = 5'h17 == _T_565 ? _next_reg_T_106 : _GEN_3428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3493 = 5'h18 == _T_565 ? _next_reg_T_106 : _GEN_3429; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3494 = 5'h19 == _T_565 ? _next_reg_T_106 : _GEN_3430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3495 = 5'h1a == _T_565 ? _next_reg_T_106 : _GEN_3431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3496 = 5'h1b == _T_565 ? _next_reg_T_106 : _GEN_3432; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3497 = 5'h1c == _T_565 ? _next_reg_T_106 : _GEN_3433; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3498 = 5'h1d == _T_565 ? _next_reg_T_106 : _GEN_3434; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3499 = 5'h1e == _T_565 ? _next_reg_T_106 : _GEN_3435; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [31:0] _GEN_3500 = 5'h1f == _T_565 ? _next_reg_T_106 : _GEN_3436; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [2:0] _GEN_3502 = _T_733 ? inst[15:13] : _GEN_3398; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3503 = _T_733 ? inst[12:10] : _GEN_3399; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3505 = _T_733 ? inst[6:2] : _GEN_3401; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3506 = _T_733 ? inst[1:0] : _GEN_3402; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3509 = _T_733 ? _GEN_3469 : _GEN_3405; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3510 = _T_733 ? _GEN_3470 : _GEN_3406; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3511 = _T_733 ? _GEN_3471 : _GEN_3407; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3512 = _T_733 ? _GEN_3472 : _GEN_3408; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3513 = _T_733 ? _GEN_3473 : _GEN_3409; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3514 = _T_733 ? _GEN_3474 : _GEN_3410; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3515 = _T_733 ? _GEN_3475 : _GEN_3411; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3516 = _T_733 ? _GEN_3476 : _GEN_3412; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3517 = _T_733 ? _GEN_3477 : _GEN_3413; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3518 = _T_733 ? _GEN_3478 : _GEN_3414; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3519 = _T_733 ? _GEN_3479 : _GEN_3415; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3520 = _T_733 ? _GEN_3480 : _GEN_3416; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3521 = _T_733 ? _GEN_3481 : _GEN_3417; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3522 = _T_733 ? _GEN_3482 : _GEN_3418; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3523 = _T_733 ? _GEN_3483 : _GEN_3419; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3524 = _T_733 ? _GEN_3484 : _GEN_3420; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3525 = _T_733 ? _GEN_3485 : _GEN_3421; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3526 = _T_733 ? _GEN_3486 : _GEN_3422; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3527 = _T_733 ? _GEN_3487 : _GEN_3423; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3528 = _T_733 ? _GEN_3488 : _GEN_3424; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3529 = _T_733 ? _GEN_3489 : _GEN_3425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3530 = _T_733 ? _GEN_3490 : _GEN_3426; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3531 = _T_733 ? _GEN_3491 : _GEN_3427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3532 = _T_733 ? _GEN_3492 : _GEN_3428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3533 = _T_733 ? _GEN_3493 : _GEN_3429; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3534 = _T_733 ? _GEN_3494 : _GEN_3430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3535 = _T_733 ? _GEN_3495 : _GEN_3431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3536 = _T_733 ? _GEN_3496 : _GEN_3432; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3537 = _T_733 ? _GEN_3497 : _GEN_3433; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3538 = _T_733 ? _GEN_3498 : _GEN_3434; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3539 = _T_733 ? _GEN_3499 : _GEN_3435; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [31:0] _GEN_3540 = _T_733 ? _GEN_3500 : _GEN_3436; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [2:0] _funct3_T_53 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _ph3_T_6 = inst[12:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_745 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_10 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_746 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_747 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_107 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_3541 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3542 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3543 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3544 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3545 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3546 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3547 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3548 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3549 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3550 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3551 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3552 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3553 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3554 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3555 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3556 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3557 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3558 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3559 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3560 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3561 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3562 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3563 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3564 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3565 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3566 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3567 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3568 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3569 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3570 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3571 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _GEN_3572 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _now_reg_next_reg_T_107 = _GEN_3364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{51,51}]
  wire [31:0] _next_reg_T_108 = _GEN_3364 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:51]
  wire [31:0] _next_reg_T_747 = _GEN_3364 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:51]
  wire [31:0] _GEN_3573 = 5'h0 == _T_565 ? _next_reg_T_108 : _GEN_3509; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3574 = 5'h1 == _T_565 ? _next_reg_T_108 : _GEN_3510; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3575 = 5'h2 == _T_565 ? _next_reg_T_108 : _GEN_3511; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3576 = 5'h3 == _T_565 ? _next_reg_T_108 : _GEN_3512; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3577 = 5'h4 == _T_565 ? _next_reg_T_108 : _GEN_3513; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3578 = 5'h5 == _T_565 ? _next_reg_T_108 : _GEN_3514; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3579 = 5'h6 == _T_565 ? _next_reg_T_108 : _GEN_3515; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3580 = 5'h7 == _T_565 ? _next_reg_T_108 : _GEN_3516; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3581 = 5'h8 == _T_565 ? _next_reg_T_108 : _GEN_3517; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3582 = 5'h9 == _T_565 ? _next_reg_T_108 : _GEN_3518; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3583 = 5'ha == _T_565 ? _next_reg_T_108 : _GEN_3519; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3584 = 5'hb == _T_565 ? _next_reg_T_108 : _GEN_3520; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3585 = 5'hc == _T_565 ? _next_reg_T_108 : _GEN_3521; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3586 = 5'hd == _T_565 ? _next_reg_T_108 : _GEN_3522; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3587 = 5'he == _T_565 ? _next_reg_T_108 : _GEN_3523; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3588 = 5'hf == _T_565 ? _next_reg_T_108 : _GEN_3524; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3589 = 5'h10 == _T_565 ? _next_reg_T_108 : _GEN_3525; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3590 = 5'h11 == _T_565 ? _next_reg_T_108 : _GEN_3526; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3591 = 5'h12 == _T_565 ? _next_reg_T_108 : _GEN_3527; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3592 = 5'h13 == _T_565 ? _next_reg_T_108 : _GEN_3528; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3593 = 5'h14 == _T_565 ? _next_reg_T_108 : _GEN_3529; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3594 = 5'h15 == _T_565 ? _next_reg_T_108 : _GEN_3530; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3595 = 5'h16 == _T_565 ? _next_reg_T_108 : _GEN_3531; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3596 = 5'h17 == _T_565 ? _next_reg_T_108 : _GEN_3532; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3597 = 5'h18 == _T_565 ? _next_reg_T_108 : _GEN_3533; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3598 = 5'h19 == _T_565 ? _next_reg_T_108 : _GEN_3534; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3599 = 5'h1a == _T_565 ? _next_reg_T_108 : _GEN_3535; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3600 = 5'h1b == _T_565 ? _next_reg_T_108 : _GEN_3536; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3601 = 5'h1c == _T_565 ? _next_reg_T_108 : _GEN_3537; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3602 = 5'h1d == _T_565 ? _next_reg_T_108 : _GEN_3538; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3603 = 5'h1e == _T_565 ? _next_reg_T_108 : _GEN_3539; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [31:0] _GEN_3604 = 5'h1f == _T_565 ? _next_reg_T_108 : _GEN_3540; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [2:0] _GEN_3606 = _T_741 ? inst[15:13] : _GEN_3502; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3607 = _T_741 ? inst[12:10] : _GEN_3503; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3609 = _T_741 ? inst[6:2] : _GEN_3505; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3610 = _T_741 ? inst[1:0] : _GEN_3506; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3613 = _T_741 ? _GEN_3573 : _GEN_3509; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3614 = _T_741 ? _GEN_3574 : _GEN_3510; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3615 = _T_741 ? _GEN_3575 : _GEN_3511; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3616 = _T_741 ? _GEN_3576 : _GEN_3512; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3617 = _T_741 ? _GEN_3577 : _GEN_3513; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3618 = _T_741 ? _GEN_3578 : _GEN_3514; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3619 = _T_741 ? _GEN_3579 : _GEN_3515; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3620 = _T_741 ? _GEN_3580 : _GEN_3516; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3621 = _T_741 ? _GEN_3581 : _GEN_3517; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3622 = _T_741 ? _GEN_3582 : _GEN_3518; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3623 = _T_741 ? _GEN_3583 : _GEN_3519; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3624 = _T_741 ? _GEN_3584 : _GEN_3520; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3625 = _T_741 ? _GEN_3585 : _GEN_3521; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3626 = _T_741 ? _GEN_3586 : _GEN_3522; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3627 = _T_741 ? _GEN_3587 : _GEN_3523; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3628 = _T_741 ? _GEN_3588 : _GEN_3524; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3629 = _T_741 ? _GEN_3589 : _GEN_3525; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3630 = _T_741 ? _GEN_3590 : _GEN_3526; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3631 = _T_741 ? _GEN_3591 : _GEN_3527; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3632 = _T_741 ? _GEN_3592 : _GEN_3528; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3633 = _T_741 ? _GEN_3593 : _GEN_3529; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3634 = _T_741 ? _GEN_3594 : _GEN_3530; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3635 = _T_741 ? _GEN_3595 : _GEN_3531; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3636 = _T_741 ? _GEN_3596 : _GEN_3532; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3637 = _T_741 ? _GEN_3597 : _GEN_3533; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3638 = _T_741 ? _GEN_3598 : _GEN_3534; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3639 = _T_741 ? _GEN_3599 : _GEN_3535; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3640 = _T_741 ? _GEN_3600 : _GEN_3536; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3641 = _T_741 ? _GEN_3601 : _GEN_3537; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3642 = _T_741 ? _GEN_3602 : _GEN_3538; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3643 = _T_741 ? _GEN_3603 : _GEN_3539; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [31:0] _GEN_3644 = _T_741 ? _GEN_3604 : _GEN_3540; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [3:0] _funct4_T_2 = inst[15:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_759 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs2_19 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_109 = io_now_reg_0 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:64]
  wire [31:0] _next_reg_T_110 = io_now_reg_0 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:64]
  wire [31:0] _next_reg_rd_32 = io_now_reg_0 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:64]
  wire [31:0] _GEN_3645 = 5'h0 == rd ? _next_reg_T_110 : _GEN_3613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3646 = 5'h1 == rd ? _next_reg_T_110 : _GEN_3614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3647 = 5'h2 == rd ? _next_reg_T_110 : _GEN_3615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3648 = 5'h3 == rd ? _next_reg_T_110 : _GEN_3616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3649 = 5'h4 == rd ? _next_reg_T_110 : _GEN_3617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3650 = 5'h5 == rd ? _next_reg_T_110 : _GEN_3618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3651 = 5'h6 == rd ? _next_reg_T_110 : _GEN_3619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3652 = 5'h7 == rd ? _next_reg_T_110 : _GEN_3620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3653 = 5'h8 == rd ? _next_reg_T_110 : _GEN_3621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3654 = 5'h9 == rd ? _next_reg_T_110 : _GEN_3622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3655 = 5'ha == rd ? _next_reg_T_110 : _GEN_3623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3656 = 5'hb == rd ? _next_reg_T_110 : _GEN_3624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3657 = 5'hc == rd ? _next_reg_T_110 : _GEN_3625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3658 = 5'hd == rd ? _next_reg_T_110 : _GEN_3626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3659 = 5'he == rd ? _next_reg_T_110 : _GEN_3627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3660 = 5'hf == rd ? _next_reg_T_110 : _GEN_3628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3661 = 5'h10 == rd ? _next_reg_T_110 : _GEN_3629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3662 = 5'h11 == rd ? _next_reg_T_110 : _GEN_3630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3663 = 5'h12 == rd ? _next_reg_T_110 : _GEN_3631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3664 = 5'h13 == rd ? _next_reg_T_110 : _GEN_3632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3665 = 5'h14 == rd ? _next_reg_T_110 : _GEN_3633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3666 = 5'h15 == rd ? _next_reg_T_110 : _GEN_3634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3667 = 5'h16 == rd ? _next_reg_T_110 : _GEN_3635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3668 = 5'h17 == rd ? _next_reg_T_110 : _GEN_3636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3669 = 5'h18 == rd ? _next_reg_T_110 : _GEN_3637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3670 = 5'h19 == rd ? _next_reg_T_110 : _GEN_3638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3671 = 5'h1a == rd ? _next_reg_T_110 : _GEN_3639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3672 = 5'h1b == rd ? _next_reg_T_110 : _GEN_3640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3673 = 5'h1c == rd ? _next_reg_T_110 : _GEN_3641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3674 = 5'h1d == rd ? _next_reg_T_110 : _GEN_3642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3675 = 5'h1e == rd ? _next_reg_T_110 : _GEN_3643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [31:0] _GEN_3676 = 5'h1f == rd ? _next_reg_T_110 : _GEN_3644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [3:0] _GEN_3678 = _T_755 ? inst[15:12] : _GEN_2842; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3681 = _T_755 ? inst[1:0] : _GEN_3610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3683 = _T_755 ? _GEN_3645 : _GEN_3613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3684 = _T_755 ? _GEN_3646 : _GEN_3614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3685 = _T_755 ? _GEN_3647 : _GEN_3615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3686 = _T_755 ? _GEN_3648 : _GEN_3616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3687 = _T_755 ? _GEN_3649 : _GEN_3617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3688 = _T_755 ? _GEN_3650 : _GEN_3618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3689 = _T_755 ? _GEN_3651 : _GEN_3619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3690 = _T_755 ? _GEN_3652 : _GEN_3620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3691 = _T_755 ? _GEN_3653 : _GEN_3621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3692 = _T_755 ? _GEN_3654 : _GEN_3622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3693 = _T_755 ? _GEN_3655 : _GEN_3623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3694 = _T_755 ? _GEN_3656 : _GEN_3624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3695 = _T_755 ? _GEN_3657 : _GEN_3625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3696 = _T_755 ? _GEN_3658 : _GEN_3626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3697 = _T_755 ? _GEN_3659 : _GEN_3627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3698 = _T_755 ? _GEN_3660 : _GEN_3628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3699 = _T_755 ? _GEN_3661 : _GEN_3629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3700 = _T_755 ? _GEN_3662 : _GEN_3630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3701 = _T_755 ? _GEN_3663 : _GEN_3631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3702 = _T_755 ? _GEN_3664 : _GEN_3632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3703 = _T_755 ? _GEN_3665 : _GEN_3633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3704 = _T_755 ? _GEN_3666 : _GEN_3634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3705 = _T_755 ? _GEN_3667 : _GEN_3635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3706 = _T_755 ? _GEN_3668 : _GEN_3636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3707 = _T_755 ? _GEN_3669 : _GEN_3637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3708 = _T_755 ? _GEN_3670 : _GEN_3638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3709 = _T_755 ? _GEN_3671 : _GEN_3639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3710 = _T_755 ? _GEN_3672 : _GEN_3640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3711 = _T_755 ? _GEN_3673 : _GEN_3641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3712 = _T_755 ? _GEN_3674 : _GEN_3642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3713 = _T_755 ? _GEN_3675 : _GEN_3643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [31:0] _GEN_3714 = _T_755 ? _GEN_3676 : _GEN_3644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [3:0] _funct4_T_3 = inst[15:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_771 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rd_1 = 5'h1f == rd ? io_now_reg_31 : _GEN_3111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [31:0] _now_reg_rs2_20 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_111 = _GEN_3112 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:63]
  wire [31:0] _next_reg_T_112 = _GEN_3112 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:63]
  wire [31:0] _next_reg_rd_33 = _GEN_3112 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:63]
  wire [31:0] _GEN_3715 = 5'h0 == rd ? _next_reg_T_112 : _GEN_3683; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3716 = 5'h1 == rd ? _next_reg_T_112 : _GEN_3684; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3717 = 5'h2 == rd ? _next_reg_T_112 : _GEN_3685; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3718 = 5'h3 == rd ? _next_reg_T_112 : _GEN_3686; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3719 = 5'h4 == rd ? _next_reg_T_112 : _GEN_3687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3720 = 5'h5 == rd ? _next_reg_T_112 : _GEN_3688; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3721 = 5'h6 == rd ? _next_reg_T_112 : _GEN_3689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3722 = 5'h7 == rd ? _next_reg_T_112 : _GEN_3690; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3723 = 5'h8 == rd ? _next_reg_T_112 : _GEN_3691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3724 = 5'h9 == rd ? _next_reg_T_112 : _GEN_3692; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3725 = 5'ha == rd ? _next_reg_T_112 : _GEN_3693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3726 = 5'hb == rd ? _next_reg_T_112 : _GEN_3694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3727 = 5'hc == rd ? _next_reg_T_112 : _GEN_3695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3728 = 5'hd == rd ? _next_reg_T_112 : _GEN_3696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3729 = 5'he == rd ? _next_reg_T_112 : _GEN_3697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3730 = 5'hf == rd ? _next_reg_T_112 : _GEN_3698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3731 = 5'h10 == rd ? _next_reg_T_112 : _GEN_3699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3732 = 5'h11 == rd ? _next_reg_T_112 : _GEN_3700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3733 = 5'h12 == rd ? _next_reg_T_112 : _GEN_3701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3734 = 5'h13 == rd ? _next_reg_T_112 : _GEN_3702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3735 = 5'h14 == rd ? _next_reg_T_112 : _GEN_3703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3736 = 5'h15 == rd ? _next_reg_T_112 : _GEN_3704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3737 = 5'h16 == rd ? _next_reg_T_112 : _GEN_3705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3738 = 5'h17 == rd ? _next_reg_T_112 : _GEN_3706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3739 = 5'h18 == rd ? _next_reg_T_112 : _GEN_3707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3740 = 5'h19 == rd ? _next_reg_T_112 : _GEN_3708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3741 = 5'h1a == rd ? _next_reg_T_112 : _GEN_3709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3742 = 5'h1b == rd ? _next_reg_T_112 : _GEN_3710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3743 = 5'h1c == rd ? _next_reg_T_112 : _GEN_3711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3744 = 5'h1d == rd ? _next_reg_T_112 : _GEN_3712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3745 = 5'h1e == rd ? _next_reg_T_112 : _GEN_3713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [31:0] _GEN_3746 = 5'h1f == rd ? _next_reg_T_112 : _GEN_3714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [3:0] _GEN_3748 = _T_767 ? inst[15:12] : _GEN_3678; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_3751 = _T_767 ? inst[1:0] : _GEN_3681; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3753 = _T_767 ? _GEN_3715 : _GEN_3683; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3754 = _T_767 ? _GEN_3716 : _GEN_3684; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3755 = _T_767 ? _GEN_3717 : _GEN_3685; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3756 = _T_767 ? _GEN_3718 : _GEN_3686; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3757 = _T_767 ? _GEN_3719 : _GEN_3687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3758 = _T_767 ? _GEN_3720 : _GEN_3688; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3759 = _T_767 ? _GEN_3721 : _GEN_3689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3760 = _T_767 ? _GEN_3722 : _GEN_3690; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3761 = _T_767 ? _GEN_3723 : _GEN_3691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3762 = _T_767 ? _GEN_3724 : _GEN_3692; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3763 = _T_767 ? _GEN_3725 : _GEN_3693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3764 = _T_767 ? _GEN_3726 : _GEN_3694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3765 = _T_767 ? _GEN_3727 : _GEN_3695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3766 = _T_767 ? _GEN_3728 : _GEN_3696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3767 = _T_767 ? _GEN_3729 : _GEN_3697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3768 = _T_767 ? _GEN_3730 : _GEN_3698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3769 = _T_767 ? _GEN_3731 : _GEN_3699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3770 = _T_767 ? _GEN_3732 : _GEN_3700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3771 = _T_767 ? _GEN_3733 : _GEN_3701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3772 = _T_767 ? _GEN_3734 : _GEN_3702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3773 = _T_767 ? _GEN_3735 : _GEN_3703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3774 = _T_767 ? _GEN_3736 : _GEN_3704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3775 = _T_767 ? _GEN_3737 : _GEN_3705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3776 = _T_767 ? _GEN_3738 : _GEN_3706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3777 = _T_767 ? _GEN_3739 : _GEN_3707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3778 = _T_767 ? _GEN_3740 : _GEN_3708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3779 = _T_767 ? _GEN_3741 : _GEN_3709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3780 = _T_767 ? _GEN_3742 : _GEN_3710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3781 = _T_767 ? _GEN_3743 : _GEN_3711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3782 = _T_767 ? _GEN_3744 : _GEN_3712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3783 = _T_767 ? _GEN_3745 : _GEN_3713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [31:0] _GEN_3784 = _T_767 ? _GEN_3746 : _GEN_3714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [5:0] _funct6_T = inst[15:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _funct2_T = inst[6:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_778 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_779 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_113 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_114 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_3785 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3786 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3787 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3788 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3789 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3790 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3791 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3792 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3793 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3794 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3795 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3796 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3797 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3798 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3799 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3800 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3801 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3802 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3803 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3804 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3805 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3806 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3807 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3808 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3809 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3810 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3811 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3812 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3813 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3814 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3815 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3816 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3817 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3818 = 5'h1 == _T_577 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3819 = 5'h2 == _T_577 ? io_now_reg_2 : _GEN_2775; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3820 = 5'h3 == _T_577 ? io_now_reg_3 : _GEN_2776; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3821 = 5'h4 == _T_577 ? io_now_reg_4 : _GEN_2777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3822 = 5'h5 == _T_577 ? io_now_reg_5 : _GEN_2778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3823 = 5'h6 == _T_577 ? io_now_reg_6 : _GEN_2779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3824 = 5'h7 == _T_577 ? io_now_reg_7 : _GEN_2780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3825 = 5'h8 == _T_577 ? io_now_reg_8 : _GEN_2781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3826 = 5'h9 == _T_577 ? io_now_reg_9 : _GEN_2782; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3827 = 5'ha == _T_577 ? io_now_reg_10 : _GEN_2783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3828 = 5'hb == _T_577 ? io_now_reg_11 : _GEN_2784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3829 = 5'hc == _T_577 ? io_now_reg_12 : _GEN_2785; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3830 = 5'hd == _T_577 ? io_now_reg_13 : _GEN_2786; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3831 = 5'he == _T_577 ? io_now_reg_14 : _GEN_2787; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3832 = 5'hf == _T_577 ? io_now_reg_15 : _GEN_2788; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3833 = 5'h10 == _T_577 ? io_now_reg_16 : _GEN_2789; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3834 = 5'h11 == _T_577 ? io_now_reg_17 : _GEN_2790; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3835 = 5'h12 == _T_577 ? io_now_reg_18 : _GEN_2791; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3836 = 5'h13 == _T_577 ? io_now_reg_19 : _GEN_2792; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3837 = 5'h14 == _T_577 ? io_now_reg_20 : _GEN_2793; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3838 = 5'h15 == _T_577 ? io_now_reg_21 : _GEN_2794; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3839 = 5'h16 == _T_577 ? io_now_reg_22 : _GEN_2795; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3840 = 5'h17 == _T_577 ? io_now_reg_23 : _GEN_2796; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3841 = 5'h18 == _T_577 ? io_now_reg_24 : _GEN_2797; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3842 = 5'h19 == _T_577 ? io_now_reg_25 : _GEN_2798; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3843 = 5'h1a == _T_577 ? io_now_reg_26 : _GEN_2799; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3844 = 5'h1b == _T_577 ? io_now_reg_27 : _GEN_2800; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3845 = 5'h1c == _T_577 ? io_now_reg_28 : _GEN_2801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3846 = 5'h1d == _T_577 ? io_now_reg_29 : _GEN_2802; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3847 = 5'h1e == _T_577 ? io_now_reg_30 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _GEN_3848 = 5'h1f == _T_577 ? io_now_reg_31 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _now_reg_next_reg_T_113 = _GEN_3364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _now_reg_next_reg_T_114 = _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{79,79}]
  wire [31:0] _next_reg_T_115 = _GEN_3364 & _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:79]
  wire [31:0] _next_reg_T_779 = _GEN_3364 & _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:79]
  wire [31:0] _GEN_3849 = 5'h0 == _T_565 ? _next_reg_T_115 : _GEN_3753; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3850 = 5'h1 == _T_565 ? _next_reg_T_115 : _GEN_3754; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3851 = 5'h2 == _T_565 ? _next_reg_T_115 : _GEN_3755; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3852 = 5'h3 == _T_565 ? _next_reg_T_115 : _GEN_3756; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3853 = 5'h4 == _T_565 ? _next_reg_T_115 : _GEN_3757; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3854 = 5'h5 == _T_565 ? _next_reg_T_115 : _GEN_3758; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3855 = 5'h6 == _T_565 ? _next_reg_T_115 : _GEN_3759; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3856 = 5'h7 == _T_565 ? _next_reg_T_115 : _GEN_3760; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3857 = 5'h8 == _T_565 ? _next_reg_T_115 : _GEN_3761; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3858 = 5'h9 == _T_565 ? _next_reg_T_115 : _GEN_3762; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3859 = 5'ha == _T_565 ? _next_reg_T_115 : _GEN_3763; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3860 = 5'hb == _T_565 ? _next_reg_T_115 : _GEN_3764; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3861 = 5'hc == _T_565 ? _next_reg_T_115 : _GEN_3765; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3862 = 5'hd == _T_565 ? _next_reg_T_115 : _GEN_3766; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3863 = 5'he == _T_565 ? _next_reg_T_115 : _GEN_3767; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3864 = 5'hf == _T_565 ? _next_reg_T_115 : _GEN_3768; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3865 = 5'h10 == _T_565 ? _next_reg_T_115 : _GEN_3769; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3866 = 5'h11 == _T_565 ? _next_reg_T_115 : _GEN_3770; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3867 = 5'h12 == _T_565 ? _next_reg_T_115 : _GEN_3771; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3868 = 5'h13 == _T_565 ? _next_reg_T_115 : _GEN_3772; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3869 = 5'h14 == _T_565 ? _next_reg_T_115 : _GEN_3773; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3870 = 5'h15 == _T_565 ? _next_reg_T_115 : _GEN_3774; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3871 = 5'h16 == _T_565 ? _next_reg_T_115 : _GEN_3775; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3872 = 5'h17 == _T_565 ? _next_reg_T_115 : _GEN_3776; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3873 = 5'h18 == _T_565 ? _next_reg_T_115 : _GEN_3777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3874 = 5'h19 == _T_565 ? _next_reg_T_115 : _GEN_3778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3875 = 5'h1a == _T_565 ? _next_reg_T_115 : _GEN_3779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3876 = 5'h1b == _T_565 ? _next_reg_T_115 : _GEN_3780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3877 = 5'h1c == _T_565 ? _next_reg_T_115 : _GEN_3781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3878 = 5'h1d == _T_565 ? _next_reg_T_115 : _GEN_3782; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3879 = 5'h1e == _T_565 ? _next_reg_T_115 : _GEN_3783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [31:0] _GEN_3880 = 5'h1f == _T_565 ? _next_reg_T_115 : _GEN_3784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [5:0] _GEN_3882 = _T_773 ? inst[15:10] : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 96:24]
  wire [1:0] _GEN_3884 = _T_773 ? inst[6:5] : 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 94:24]
  wire [1:0] _GEN_3886 = _T_773 ? inst[1:0] : _GEN_3751; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3888 = _T_773 ? _GEN_3849 : _GEN_3753; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3889 = _T_773 ? _GEN_3850 : _GEN_3754; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3890 = _T_773 ? _GEN_3851 : _GEN_3755; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3891 = _T_773 ? _GEN_3852 : _GEN_3756; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3892 = _T_773 ? _GEN_3853 : _GEN_3757; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3893 = _T_773 ? _GEN_3854 : _GEN_3758; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3894 = _T_773 ? _GEN_3855 : _GEN_3759; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3895 = _T_773 ? _GEN_3856 : _GEN_3760; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3896 = _T_773 ? _GEN_3857 : _GEN_3761; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3897 = _T_773 ? _GEN_3858 : _GEN_3762; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3898 = _T_773 ? _GEN_3859 : _GEN_3763; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3899 = _T_773 ? _GEN_3860 : _GEN_3764; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3900 = _T_773 ? _GEN_3861 : _GEN_3765; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3901 = _T_773 ? _GEN_3862 : _GEN_3766; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3902 = _T_773 ? _GEN_3863 : _GEN_3767; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3903 = _T_773 ? _GEN_3864 : _GEN_3768; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3904 = _T_773 ? _GEN_3865 : _GEN_3769; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3905 = _T_773 ? _GEN_3866 : _GEN_3770; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3906 = _T_773 ? _GEN_3867 : _GEN_3771; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3907 = _T_773 ? _GEN_3868 : _GEN_3772; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3908 = _T_773 ? _GEN_3869 : _GEN_3773; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3909 = _T_773 ? _GEN_3870 : _GEN_3774; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3910 = _T_773 ? _GEN_3871 : _GEN_3775; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3911 = _T_773 ? _GEN_3872 : _GEN_3776; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3912 = _T_773 ? _GEN_3873 : _GEN_3777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3913 = _T_773 ? _GEN_3874 : _GEN_3778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3914 = _T_773 ? _GEN_3875 : _GEN_3779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3915 = _T_773 ? _GEN_3876 : _GEN_3780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3916 = _T_773 ? _GEN_3877 : _GEN_3781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3917 = _T_773 ? _GEN_3878 : _GEN_3782; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3918 = _T_773 ? _GEN_3879 : _GEN_3783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [31:0] _GEN_3919 = _T_773 ? _GEN_3880 : _GEN_3784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [5:0] _funct6_T_1 = inst[15:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _funct2_T_1 = inst[6:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_786 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_787 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_116 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_117 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_3920 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3921 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3922 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3923 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3924 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3925 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3926 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3927 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3928 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3929 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3930 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3931 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3932 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3933 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3934 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3935 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3936 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3937 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3938 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3939 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3940 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3941 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3942 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3943 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3944 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3945 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3946 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3947 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3948 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3949 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3950 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3951 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3952 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3953 = 5'h1 == _T_577 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3954 = 5'h2 == _T_577 ? io_now_reg_2 : _GEN_2775; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3955 = 5'h3 == _T_577 ? io_now_reg_3 : _GEN_2776; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3956 = 5'h4 == _T_577 ? io_now_reg_4 : _GEN_2777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3957 = 5'h5 == _T_577 ? io_now_reg_5 : _GEN_2778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3958 = 5'h6 == _T_577 ? io_now_reg_6 : _GEN_2779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3959 = 5'h7 == _T_577 ? io_now_reg_7 : _GEN_2780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3960 = 5'h8 == _T_577 ? io_now_reg_8 : _GEN_2781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3961 = 5'h9 == _T_577 ? io_now_reg_9 : _GEN_2782; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3962 = 5'ha == _T_577 ? io_now_reg_10 : _GEN_2783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3963 = 5'hb == _T_577 ? io_now_reg_11 : _GEN_2784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3964 = 5'hc == _T_577 ? io_now_reg_12 : _GEN_2785; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3965 = 5'hd == _T_577 ? io_now_reg_13 : _GEN_2786; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3966 = 5'he == _T_577 ? io_now_reg_14 : _GEN_2787; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3967 = 5'hf == _T_577 ? io_now_reg_15 : _GEN_2788; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3968 = 5'h10 == _T_577 ? io_now_reg_16 : _GEN_2789; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3969 = 5'h11 == _T_577 ? io_now_reg_17 : _GEN_2790; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3970 = 5'h12 == _T_577 ? io_now_reg_18 : _GEN_2791; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3971 = 5'h13 == _T_577 ? io_now_reg_19 : _GEN_2792; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3972 = 5'h14 == _T_577 ? io_now_reg_20 : _GEN_2793; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3973 = 5'h15 == _T_577 ? io_now_reg_21 : _GEN_2794; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3974 = 5'h16 == _T_577 ? io_now_reg_22 : _GEN_2795; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3975 = 5'h17 == _T_577 ? io_now_reg_23 : _GEN_2796; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3976 = 5'h18 == _T_577 ? io_now_reg_24 : _GEN_2797; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3977 = 5'h19 == _T_577 ? io_now_reg_25 : _GEN_2798; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3978 = 5'h1a == _T_577 ? io_now_reg_26 : _GEN_2799; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3979 = 5'h1b == _T_577 ? io_now_reg_27 : _GEN_2800; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3980 = 5'h1c == _T_577 ? io_now_reg_28 : _GEN_2801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3981 = 5'h1d == _T_577 ? io_now_reg_29 : _GEN_2802; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3982 = 5'h1e == _T_577 ? io_now_reg_30 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _GEN_3983 = 5'h1f == _T_577 ? io_now_reg_31 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _now_reg_next_reg_T_116 = _GEN_3364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _now_reg_next_reg_T_117 = _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{79,79}]
  wire [31:0] _next_reg_T_118 = _GEN_3364 | _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:79]
  wire [31:0] _next_reg_T_787 = _GEN_3364 | _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:79]
  wire [31:0] _GEN_3984 = 5'h0 == _T_565 ? _next_reg_T_118 : _GEN_3888; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3985 = 5'h1 == _T_565 ? _next_reg_T_118 : _GEN_3889; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3986 = 5'h2 == _T_565 ? _next_reg_T_118 : _GEN_3890; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3987 = 5'h3 == _T_565 ? _next_reg_T_118 : _GEN_3891; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3988 = 5'h4 == _T_565 ? _next_reg_T_118 : _GEN_3892; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3989 = 5'h5 == _T_565 ? _next_reg_T_118 : _GEN_3893; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3990 = 5'h6 == _T_565 ? _next_reg_T_118 : _GEN_3894; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3991 = 5'h7 == _T_565 ? _next_reg_T_118 : _GEN_3895; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3992 = 5'h8 == _T_565 ? _next_reg_T_118 : _GEN_3896; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3993 = 5'h9 == _T_565 ? _next_reg_T_118 : _GEN_3897; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3994 = 5'ha == _T_565 ? _next_reg_T_118 : _GEN_3898; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3995 = 5'hb == _T_565 ? _next_reg_T_118 : _GEN_3899; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3996 = 5'hc == _T_565 ? _next_reg_T_118 : _GEN_3900; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3997 = 5'hd == _T_565 ? _next_reg_T_118 : _GEN_3901; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3998 = 5'he == _T_565 ? _next_reg_T_118 : _GEN_3902; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_3999 = 5'hf == _T_565 ? _next_reg_T_118 : _GEN_3903; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4000 = 5'h10 == _T_565 ? _next_reg_T_118 : _GEN_3904; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4001 = 5'h11 == _T_565 ? _next_reg_T_118 : _GEN_3905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4002 = 5'h12 == _T_565 ? _next_reg_T_118 : _GEN_3906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4003 = 5'h13 == _T_565 ? _next_reg_T_118 : _GEN_3907; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4004 = 5'h14 == _T_565 ? _next_reg_T_118 : _GEN_3908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4005 = 5'h15 == _T_565 ? _next_reg_T_118 : _GEN_3909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4006 = 5'h16 == _T_565 ? _next_reg_T_118 : _GEN_3910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4007 = 5'h17 == _T_565 ? _next_reg_T_118 : _GEN_3911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4008 = 5'h18 == _T_565 ? _next_reg_T_118 : _GEN_3912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4009 = 5'h19 == _T_565 ? _next_reg_T_118 : _GEN_3913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4010 = 5'h1a == _T_565 ? _next_reg_T_118 : _GEN_3914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4011 = 5'h1b == _T_565 ? _next_reg_T_118 : _GEN_3915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4012 = 5'h1c == _T_565 ? _next_reg_T_118 : _GEN_3916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4013 = 5'h1d == _T_565 ? _next_reg_T_118 : _GEN_3917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4014 = 5'h1e == _T_565 ? _next_reg_T_118 : _GEN_3918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [31:0] _GEN_4015 = 5'h1f == _T_565 ? _next_reg_T_118 : _GEN_3919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [5:0] _GEN_4017 = _T_781 ? inst[15:10] : _GEN_3882; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4019 = _T_781 ? inst[6:5] : _GEN_3884; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4021 = _T_781 ? inst[1:0] : _GEN_3886; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4023 = _T_781 ? _GEN_3984 : _GEN_3888; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4024 = _T_781 ? _GEN_3985 : _GEN_3889; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4025 = _T_781 ? _GEN_3986 : _GEN_3890; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4026 = _T_781 ? _GEN_3987 : _GEN_3891; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4027 = _T_781 ? _GEN_3988 : _GEN_3892; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4028 = _T_781 ? _GEN_3989 : _GEN_3893; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4029 = _T_781 ? _GEN_3990 : _GEN_3894; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4030 = _T_781 ? _GEN_3991 : _GEN_3895; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4031 = _T_781 ? _GEN_3992 : _GEN_3896; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4032 = _T_781 ? _GEN_3993 : _GEN_3897; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4033 = _T_781 ? _GEN_3994 : _GEN_3898; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4034 = _T_781 ? _GEN_3995 : _GEN_3899; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4035 = _T_781 ? _GEN_3996 : _GEN_3900; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4036 = _T_781 ? _GEN_3997 : _GEN_3901; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4037 = _T_781 ? _GEN_3998 : _GEN_3902; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4038 = _T_781 ? _GEN_3999 : _GEN_3903; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4039 = _T_781 ? _GEN_4000 : _GEN_3904; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4040 = _T_781 ? _GEN_4001 : _GEN_3905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4041 = _T_781 ? _GEN_4002 : _GEN_3906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4042 = _T_781 ? _GEN_4003 : _GEN_3907; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4043 = _T_781 ? _GEN_4004 : _GEN_3908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4044 = _T_781 ? _GEN_4005 : _GEN_3909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4045 = _T_781 ? _GEN_4006 : _GEN_3910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4046 = _T_781 ? _GEN_4007 : _GEN_3911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4047 = _T_781 ? _GEN_4008 : _GEN_3912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4048 = _T_781 ? _GEN_4009 : _GEN_3913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4049 = _T_781 ? _GEN_4010 : _GEN_3914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4050 = _T_781 ? _GEN_4011 : _GEN_3915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4051 = _T_781 ? _GEN_4012 : _GEN_3916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4052 = _T_781 ? _GEN_4013 : _GEN_3917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4053 = _T_781 ? _GEN_4014 : _GEN_3918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [31:0] _GEN_4054 = _T_781 ? _GEN_4015 : _GEN_3919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [5:0] _funct6_T_2 = inst[15:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _funct2_T_2 = inst[6:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_794 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_795 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_119 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_120 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_4055 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_4056 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4057 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4058 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4059 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4060 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4061 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4062 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4063 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4064 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4065 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4066 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4067 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4068 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4069 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4070 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4071 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4072 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4073 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4074 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4075 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4076 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4077 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4078 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4079 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4080 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4081 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4082 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4083 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4084 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4085 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4086 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4087 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_4088 = 5'h1 == _T_577 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4089 = 5'h2 == _T_577 ? io_now_reg_2 : _GEN_2775; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4090 = 5'h3 == _T_577 ? io_now_reg_3 : _GEN_2776; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4091 = 5'h4 == _T_577 ? io_now_reg_4 : _GEN_2777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4092 = 5'h5 == _T_577 ? io_now_reg_5 : _GEN_2778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4093 = 5'h6 == _T_577 ? io_now_reg_6 : _GEN_2779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4094 = 5'h7 == _T_577 ? io_now_reg_7 : _GEN_2780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4095 = 5'h8 == _T_577 ? io_now_reg_8 : _GEN_2781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4096 = 5'h9 == _T_577 ? io_now_reg_9 : _GEN_2782; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4097 = 5'ha == _T_577 ? io_now_reg_10 : _GEN_2783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4098 = 5'hb == _T_577 ? io_now_reg_11 : _GEN_2784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4099 = 5'hc == _T_577 ? io_now_reg_12 : _GEN_2785; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4100 = 5'hd == _T_577 ? io_now_reg_13 : _GEN_2786; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4101 = 5'he == _T_577 ? io_now_reg_14 : _GEN_2787; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4102 = 5'hf == _T_577 ? io_now_reg_15 : _GEN_2788; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4103 = 5'h10 == _T_577 ? io_now_reg_16 : _GEN_2789; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4104 = 5'h11 == _T_577 ? io_now_reg_17 : _GEN_2790; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4105 = 5'h12 == _T_577 ? io_now_reg_18 : _GEN_2791; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4106 = 5'h13 == _T_577 ? io_now_reg_19 : _GEN_2792; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4107 = 5'h14 == _T_577 ? io_now_reg_20 : _GEN_2793; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4108 = 5'h15 == _T_577 ? io_now_reg_21 : _GEN_2794; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4109 = 5'h16 == _T_577 ? io_now_reg_22 : _GEN_2795; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4110 = 5'h17 == _T_577 ? io_now_reg_23 : _GEN_2796; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4111 = 5'h18 == _T_577 ? io_now_reg_24 : _GEN_2797; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4112 = 5'h19 == _T_577 ? io_now_reg_25 : _GEN_2798; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4113 = 5'h1a == _T_577 ? io_now_reg_26 : _GEN_2799; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4114 = 5'h1b == _T_577 ? io_now_reg_27 : _GEN_2800; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4115 = 5'h1c == _T_577 ? io_now_reg_28 : _GEN_2801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4116 = 5'h1d == _T_577 ? io_now_reg_29 : _GEN_2802; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4117 = 5'h1e == _T_577 ? io_now_reg_30 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _GEN_4118 = 5'h1f == _T_577 ? io_now_reg_31 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _now_reg_next_reg_T_119 = _GEN_3364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _now_reg_next_reg_T_120 = _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{79,79}]
  wire [31:0] _next_reg_T_121 = _GEN_3364 ^ _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:79]
  wire [31:0] _next_reg_T_795 = _GEN_3364 ^ _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:79]
  wire [31:0] _GEN_4119 = 5'h0 == _T_565 ? _next_reg_T_121 : _GEN_4023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4120 = 5'h1 == _T_565 ? _next_reg_T_121 : _GEN_4024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4121 = 5'h2 == _T_565 ? _next_reg_T_121 : _GEN_4025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4122 = 5'h3 == _T_565 ? _next_reg_T_121 : _GEN_4026; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4123 = 5'h4 == _T_565 ? _next_reg_T_121 : _GEN_4027; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4124 = 5'h5 == _T_565 ? _next_reg_T_121 : _GEN_4028; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4125 = 5'h6 == _T_565 ? _next_reg_T_121 : _GEN_4029; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4126 = 5'h7 == _T_565 ? _next_reg_T_121 : _GEN_4030; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4127 = 5'h8 == _T_565 ? _next_reg_T_121 : _GEN_4031; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4128 = 5'h9 == _T_565 ? _next_reg_T_121 : _GEN_4032; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4129 = 5'ha == _T_565 ? _next_reg_T_121 : _GEN_4033; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4130 = 5'hb == _T_565 ? _next_reg_T_121 : _GEN_4034; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4131 = 5'hc == _T_565 ? _next_reg_T_121 : _GEN_4035; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4132 = 5'hd == _T_565 ? _next_reg_T_121 : _GEN_4036; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4133 = 5'he == _T_565 ? _next_reg_T_121 : _GEN_4037; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4134 = 5'hf == _T_565 ? _next_reg_T_121 : _GEN_4038; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4135 = 5'h10 == _T_565 ? _next_reg_T_121 : _GEN_4039; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4136 = 5'h11 == _T_565 ? _next_reg_T_121 : _GEN_4040; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4137 = 5'h12 == _T_565 ? _next_reg_T_121 : _GEN_4041; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4138 = 5'h13 == _T_565 ? _next_reg_T_121 : _GEN_4042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4139 = 5'h14 == _T_565 ? _next_reg_T_121 : _GEN_4043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4140 = 5'h15 == _T_565 ? _next_reg_T_121 : _GEN_4044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4141 = 5'h16 == _T_565 ? _next_reg_T_121 : _GEN_4045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4142 = 5'h17 == _T_565 ? _next_reg_T_121 : _GEN_4046; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4143 = 5'h18 == _T_565 ? _next_reg_T_121 : _GEN_4047; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4144 = 5'h19 == _T_565 ? _next_reg_T_121 : _GEN_4048; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4145 = 5'h1a == _T_565 ? _next_reg_T_121 : _GEN_4049; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4146 = 5'h1b == _T_565 ? _next_reg_T_121 : _GEN_4050; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4147 = 5'h1c == _T_565 ? _next_reg_T_121 : _GEN_4051; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4148 = 5'h1d == _T_565 ? _next_reg_T_121 : _GEN_4052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4149 = 5'h1e == _T_565 ? _next_reg_T_121 : _GEN_4053; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [31:0] _GEN_4150 = 5'h1f == _T_565 ? _next_reg_T_121 : _GEN_4054; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [5:0] _GEN_4152 = _T_789 ? inst[15:10] : _GEN_4017; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4154 = _T_789 ? inst[6:5] : _GEN_4019; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4156 = _T_789 ? inst[1:0] : _GEN_4021; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4158 = _T_789 ? _GEN_4119 : _GEN_4023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4159 = _T_789 ? _GEN_4120 : _GEN_4024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4160 = _T_789 ? _GEN_4121 : _GEN_4025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4161 = _T_789 ? _GEN_4122 : _GEN_4026; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4162 = _T_789 ? _GEN_4123 : _GEN_4027; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4163 = _T_789 ? _GEN_4124 : _GEN_4028; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4164 = _T_789 ? _GEN_4125 : _GEN_4029; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4165 = _T_789 ? _GEN_4126 : _GEN_4030; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4166 = _T_789 ? _GEN_4127 : _GEN_4031; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4167 = _T_789 ? _GEN_4128 : _GEN_4032; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4168 = _T_789 ? _GEN_4129 : _GEN_4033; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4169 = _T_789 ? _GEN_4130 : _GEN_4034; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4170 = _T_789 ? _GEN_4131 : _GEN_4035; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4171 = _T_789 ? _GEN_4132 : _GEN_4036; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4172 = _T_789 ? _GEN_4133 : _GEN_4037; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4173 = _T_789 ? _GEN_4134 : _GEN_4038; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4174 = _T_789 ? _GEN_4135 : _GEN_4039; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4175 = _T_789 ? _GEN_4136 : _GEN_4040; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4176 = _T_789 ? _GEN_4137 : _GEN_4041; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4177 = _T_789 ? _GEN_4138 : _GEN_4042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4178 = _T_789 ? _GEN_4139 : _GEN_4043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4179 = _T_789 ? _GEN_4140 : _GEN_4044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4180 = _T_789 ? _GEN_4141 : _GEN_4045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4181 = _T_789 ? _GEN_4142 : _GEN_4046; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4182 = _T_789 ? _GEN_4143 : _GEN_4047; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4183 = _T_789 ? _GEN_4144 : _GEN_4048; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4184 = _T_789 ? _GEN_4145 : _GEN_4049; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4185 = _T_789 ? _GEN_4146 : _GEN_4050; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4186 = _T_789 ? _GEN_4147 : _GEN_4051; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4187 = _T_789 ? _GEN_4148 : _GEN_4052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4188 = _T_789 ? _GEN_4149 : _GEN_4053; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [31:0] _GEN_4189 = _T_789 ? _GEN_4150 : _GEN_4054; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [5:0] _funct6_T_3 = inst[15:10]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _funct2_T_3 = inst[6:5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_802 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _T_803 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_122 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_123 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [31:0] _GEN_4190 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_4191 = 5'h1 == _T_565 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4192 = 5'h2 == _T_565 ? io_now_reg_2 : _GEN_3334; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4193 = 5'h3 == _T_565 ? io_now_reg_3 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4194 = 5'h4 == _T_565 ? io_now_reg_4 : _GEN_3336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4195 = 5'h5 == _T_565 ? io_now_reg_5 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4196 = 5'h6 == _T_565 ? io_now_reg_6 : _GEN_3338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4197 = 5'h7 == _T_565 ? io_now_reg_7 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4198 = 5'h8 == _T_565 ? io_now_reg_8 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4199 = 5'h9 == _T_565 ? io_now_reg_9 : _GEN_3341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4200 = 5'ha == _T_565 ? io_now_reg_10 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4201 = 5'hb == _T_565 ? io_now_reg_11 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4202 = 5'hc == _T_565 ? io_now_reg_12 : _GEN_3344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4203 = 5'hd == _T_565 ? io_now_reg_13 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4204 = 5'he == _T_565 ? io_now_reg_14 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4205 = 5'hf == _T_565 ? io_now_reg_15 : _GEN_3347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4206 = 5'h10 == _T_565 ? io_now_reg_16 : _GEN_3348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4207 = 5'h11 == _T_565 ? io_now_reg_17 : _GEN_3349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4208 = 5'h12 == _T_565 ? io_now_reg_18 : _GEN_3350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4209 = 5'h13 == _T_565 ? io_now_reg_19 : _GEN_3351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4210 = 5'h14 == _T_565 ? io_now_reg_20 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4211 = 5'h15 == _T_565 ? io_now_reg_21 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4212 = 5'h16 == _T_565 ? io_now_reg_22 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4213 = 5'h17 == _T_565 ? io_now_reg_23 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4214 = 5'h18 == _T_565 ? io_now_reg_24 : _GEN_3356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4215 = 5'h19 == _T_565 ? io_now_reg_25 : _GEN_3357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4216 = 5'h1a == _T_565 ? io_now_reg_26 : _GEN_3358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4217 = 5'h1b == _T_565 ? io_now_reg_27 : _GEN_3359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4218 = 5'h1c == _T_565 ? io_now_reg_28 : _GEN_3360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4219 = 5'h1d == _T_565 ? io_now_reg_29 : _GEN_3361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4220 = 5'h1e == _T_565 ? io_now_reg_30 : _GEN_3362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4221 = 5'h1f == _T_565 ? io_now_reg_31 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4222 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_4223 = 5'h1 == _T_577 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4224 = 5'h2 == _T_577 ? io_now_reg_2 : _GEN_2775; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4225 = 5'h3 == _T_577 ? io_now_reg_3 : _GEN_2776; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4226 = 5'h4 == _T_577 ? io_now_reg_4 : _GEN_2777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4227 = 5'h5 == _T_577 ? io_now_reg_5 : _GEN_2778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4228 = 5'h6 == _T_577 ? io_now_reg_6 : _GEN_2779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4229 = 5'h7 == _T_577 ? io_now_reg_7 : _GEN_2780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4230 = 5'h8 == _T_577 ? io_now_reg_8 : _GEN_2781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4231 = 5'h9 == _T_577 ? io_now_reg_9 : _GEN_2782; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4232 = 5'ha == _T_577 ? io_now_reg_10 : _GEN_2783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4233 = 5'hb == _T_577 ? io_now_reg_11 : _GEN_2784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4234 = 5'hc == _T_577 ? io_now_reg_12 : _GEN_2785; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4235 = 5'hd == _T_577 ? io_now_reg_13 : _GEN_2786; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4236 = 5'he == _T_577 ? io_now_reg_14 : _GEN_2787; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4237 = 5'hf == _T_577 ? io_now_reg_15 : _GEN_2788; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4238 = 5'h10 == _T_577 ? io_now_reg_16 : _GEN_2789; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4239 = 5'h11 == _T_577 ? io_now_reg_17 : _GEN_2790; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4240 = 5'h12 == _T_577 ? io_now_reg_18 : _GEN_2791; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4241 = 5'h13 == _T_577 ? io_now_reg_19 : _GEN_2792; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4242 = 5'h14 == _T_577 ? io_now_reg_20 : _GEN_2793; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4243 = 5'h15 == _T_577 ? io_now_reg_21 : _GEN_2794; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4244 = 5'h16 == _T_577 ? io_now_reg_22 : _GEN_2795; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4245 = 5'h17 == _T_577 ? io_now_reg_23 : _GEN_2796; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4246 = 5'h18 == _T_577 ? io_now_reg_24 : _GEN_2797; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4247 = 5'h19 == _T_577 ? io_now_reg_25 : _GEN_2798; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4248 = 5'h1a == _T_577 ? io_now_reg_26 : _GEN_2799; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4249 = 5'h1b == _T_577 ? io_now_reg_27 : _GEN_2800; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4250 = 5'h1c == _T_577 ? io_now_reg_28 : _GEN_2801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4251 = 5'h1d == _T_577 ? io_now_reg_29 : _GEN_2802; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4252 = 5'h1e == _T_577 ? io_now_reg_30 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _GEN_4253 = 5'h1f == _T_577 ? io_now_reg_31 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _now_reg_next_reg_T_122 = _GEN_3364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [31:0] _now_reg_next_reg_T_123 = _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{79,79}]
  wire [32:0] _next_reg_T_124 = _GEN_3364 - _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:79]
  wire [31:0] _next_reg_T_125 = _GEN_3364 - _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:79]
  wire [31:0] _next_reg_T_803 = _GEN_3364 - _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:79]
  wire [31:0] _GEN_4254 = 5'h0 == _T_565 ? _next_reg_T_125 : _GEN_4158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4255 = 5'h1 == _T_565 ? _next_reg_T_125 : _GEN_4159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4256 = 5'h2 == _T_565 ? _next_reg_T_125 : _GEN_4160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4257 = 5'h3 == _T_565 ? _next_reg_T_125 : _GEN_4161; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4258 = 5'h4 == _T_565 ? _next_reg_T_125 : _GEN_4162; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4259 = 5'h5 == _T_565 ? _next_reg_T_125 : _GEN_4163; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4260 = 5'h6 == _T_565 ? _next_reg_T_125 : _GEN_4164; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4261 = 5'h7 == _T_565 ? _next_reg_T_125 : _GEN_4165; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4262 = 5'h8 == _T_565 ? _next_reg_T_125 : _GEN_4166; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4263 = 5'h9 == _T_565 ? _next_reg_T_125 : _GEN_4167; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4264 = 5'ha == _T_565 ? _next_reg_T_125 : _GEN_4168; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4265 = 5'hb == _T_565 ? _next_reg_T_125 : _GEN_4169; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4266 = 5'hc == _T_565 ? _next_reg_T_125 : _GEN_4170; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4267 = 5'hd == _T_565 ? _next_reg_T_125 : _GEN_4171; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4268 = 5'he == _T_565 ? _next_reg_T_125 : _GEN_4172; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4269 = 5'hf == _T_565 ? _next_reg_T_125 : _GEN_4173; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4270 = 5'h10 == _T_565 ? _next_reg_T_125 : _GEN_4174; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4271 = 5'h11 == _T_565 ? _next_reg_T_125 : _GEN_4175; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4272 = 5'h12 == _T_565 ? _next_reg_T_125 : _GEN_4176; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4273 = 5'h13 == _T_565 ? _next_reg_T_125 : _GEN_4177; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4274 = 5'h14 == _T_565 ? _next_reg_T_125 : _GEN_4178; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4275 = 5'h15 == _T_565 ? _next_reg_T_125 : _GEN_4179; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4276 = 5'h16 == _T_565 ? _next_reg_T_125 : _GEN_4180; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4277 = 5'h17 == _T_565 ? _next_reg_T_125 : _GEN_4181; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4278 = 5'h18 == _T_565 ? _next_reg_T_125 : _GEN_4182; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4279 = 5'h19 == _T_565 ? _next_reg_T_125 : _GEN_4183; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4280 = 5'h1a == _T_565 ? _next_reg_T_125 : _GEN_4184; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4281 = 5'h1b == _T_565 ? _next_reg_T_125 : _GEN_4185; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4282 = 5'h1c == _T_565 ? _next_reg_T_125 : _GEN_4186; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4283 = 5'h1d == _T_565 ? _next_reg_T_125 : _GEN_4187; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4284 = 5'h1e == _T_565 ? _next_reg_T_125 : _GEN_4188; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [31:0] _GEN_4285 = 5'h1f == _T_565 ? _next_reg_T_125 : _GEN_4189; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [5:0] _GEN_4287 = _T_797 ? inst[15:10] : _GEN_4152; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4289 = _T_797 ? inst[6:5] : _GEN_4154; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4291 = _T_797 ? inst[1:0] : _GEN_4156; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4293 = _T_797 ? _GEN_4254 : _GEN_4158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4294 = _T_797 ? _GEN_4255 : _GEN_4159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4295 = _T_797 ? _GEN_4256 : _GEN_4160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4296 = _T_797 ? _GEN_4257 : _GEN_4161; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4297 = _T_797 ? _GEN_4258 : _GEN_4162; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4298 = _T_797 ? _GEN_4259 : _GEN_4163; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4299 = _T_797 ? _GEN_4260 : _GEN_4164; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4300 = _T_797 ? _GEN_4261 : _GEN_4165; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4301 = _T_797 ? _GEN_4262 : _GEN_4166; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4302 = _T_797 ? _GEN_4263 : _GEN_4167; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4303 = _T_797 ? _GEN_4264 : _GEN_4168; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4304 = _T_797 ? _GEN_4265 : _GEN_4169; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4305 = _T_797 ? _GEN_4266 : _GEN_4170; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4306 = _T_797 ? _GEN_4267 : _GEN_4171; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4307 = _T_797 ? _GEN_4268 : _GEN_4172; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4308 = _T_797 ? _GEN_4269 : _GEN_4173; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4309 = _T_797 ? _GEN_4270 : _GEN_4174; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4310 = _T_797 ? _GEN_4271 : _GEN_4175; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4311 = _T_797 ? _GEN_4272 : _GEN_4176; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4312 = _T_797 ? _GEN_4273 : _GEN_4177; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4313 = _T_797 ? _GEN_4274 : _GEN_4178; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4314 = _T_797 ? _GEN_4275 : _GEN_4179; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4315 = _T_797 ? _GEN_4276 : _GEN_4180; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4316 = _T_797 ? _GEN_4277 : _GEN_4181; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4317 = _T_797 ? _GEN_4278 : _GEN_4182; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4318 = _T_797 ? _GEN_4279 : _GEN_4183; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4319 = _T_797 ? _GEN_4280 : _GEN_4184; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4320 = _T_797 ? _GEN_4281 : _GEN_4185; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4321 = _T_797 ? _GEN_4282 : _GEN_4186; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4322 = _T_797 ? _GEN_4283 : _GEN_4187; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4323 = _T_797 ? _GEN_4284 : _GEN_4188; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [31:0] _GEN_4324 = _T_797 ? _GEN_4285 : _GEN_4189; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [2:0] _funct3_T_54 = inst[15:13]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _ph1_T_6 = inst[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_809 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _ph5_T_11 = inst[6:2]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [1:0] _T_810 = inst[1:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_4326 = _T_805 ? inst[15:13] : _GEN_3606; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_4327 = _T_805 ? inst[12] : _GEN_3295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4329 = _T_805 ? inst[6:2] : _GEN_3609; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [1:0] _GEN_4330 = _T_805 ? inst[1:0] : _GEN_4291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [6:0] _funct7_T_10 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_55 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_817 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_49 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_21 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _next_reg_T_126 = _GEN_31 * _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:65]
  wire [31:0] _next_reg_T_127 = _next_reg_T_126[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:80]
  wire [31:0] _next_reg_rd_34 = _next_reg_T_126[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:80]
  wire [31:0] _GEN_4332 = 5'h0 == rd ? _next_reg_T_126[31:0] : _GEN_4293; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4333 = 5'h1 == rd ? _next_reg_T_126[31:0] : _GEN_4294; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4334 = 5'h2 == rd ? _next_reg_T_126[31:0] : _GEN_4295; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4335 = 5'h3 == rd ? _next_reg_T_126[31:0] : _GEN_4296; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4336 = 5'h4 == rd ? _next_reg_T_126[31:0] : _GEN_4297; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4337 = 5'h5 == rd ? _next_reg_T_126[31:0] : _GEN_4298; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4338 = 5'h6 == rd ? _next_reg_T_126[31:0] : _GEN_4299; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4339 = 5'h7 == rd ? _next_reg_T_126[31:0] : _GEN_4300; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4340 = 5'h8 == rd ? _next_reg_T_126[31:0] : _GEN_4301; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4341 = 5'h9 == rd ? _next_reg_T_126[31:0] : _GEN_4302; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4342 = 5'ha == rd ? _next_reg_T_126[31:0] : _GEN_4303; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4343 = 5'hb == rd ? _next_reg_T_126[31:0] : _GEN_4304; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4344 = 5'hc == rd ? _next_reg_T_126[31:0] : _GEN_4305; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4345 = 5'hd == rd ? _next_reg_T_126[31:0] : _GEN_4306; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4346 = 5'he == rd ? _next_reg_T_126[31:0] : _GEN_4307; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4347 = 5'hf == rd ? _next_reg_T_126[31:0] : _GEN_4308; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4348 = 5'h10 == rd ? _next_reg_T_126[31:0] : _GEN_4309; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4349 = 5'h11 == rd ? _next_reg_T_126[31:0] : _GEN_4310; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4350 = 5'h12 == rd ? _next_reg_T_126[31:0] : _GEN_4311; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4351 = 5'h13 == rd ? _next_reg_T_126[31:0] : _GEN_4312; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4352 = 5'h14 == rd ? _next_reg_T_126[31:0] : _GEN_4313; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4353 = 5'h15 == rd ? _next_reg_T_126[31:0] : _GEN_4314; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4354 = 5'h16 == rd ? _next_reg_T_126[31:0] : _GEN_4315; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4355 = 5'h17 == rd ? _next_reg_T_126[31:0] : _GEN_4316; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4356 = 5'h18 == rd ? _next_reg_T_126[31:0] : _GEN_4317; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4357 = 5'h19 == rd ? _next_reg_T_126[31:0] : _GEN_4318; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4358 = 5'h1a == rd ? _next_reg_T_126[31:0] : _GEN_4319; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4359 = 5'h1b == rd ? _next_reg_T_126[31:0] : _GEN_4320; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4360 = 5'h1c == rd ? _next_reg_T_126[31:0] : _GEN_4321; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4361 = 5'h1d == rd ? _next_reg_T_126[31:0] : _GEN_4322; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4362 = 5'h1e == rd ? _next_reg_T_126[31:0] : _GEN_4323; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_4363 = 5'h1f == rd ? _next_reg_T_126[31:0] : _GEN_4324; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [6:0] _GEN_4365 = _T_812 ? inst[31:25] : _GEN_1513; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4368 = _T_812 ? inst[14:12] : _GEN_4326; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4370 = _T_812 ? inst[6:0] : _GEN_2548; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4371 = _T_812 ? _GEN_4332 : _GEN_4293; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4372 = _T_812 ? _GEN_4333 : _GEN_4294; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4373 = _T_812 ? _GEN_4334 : _GEN_4295; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4374 = _T_812 ? _GEN_4335 : _GEN_4296; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4375 = _T_812 ? _GEN_4336 : _GEN_4297; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4376 = _T_812 ? _GEN_4337 : _GEN_4298; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4377 = _T_812 ? _GEN_4338 : _GEN_4299; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4378 = _T_812 ? _GEN_4339 : _GEN_4300; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4379 = _T_812 ? _GEN_4340 : _GEN_4301; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4380 = _T_812 ? _GEN_4341 : _GEN_4302; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4381 = _T_812 ? _GEN_4342 : _GEN_4303; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4382 = _T_812 ? _GEN_4343 : _GEN_4304; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4383 = _T_812 ? _GEN_4344 : _GEN_4305; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4384 = _T_812 ? _GEN_4345 : _GEN_4306; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4385 = _T_812 ? _GEN_4346 : _GEN_4307; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4386 = _T_812 ? _GEN_4347 : _GEN_4308; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4387 = _T_812 ? _GEN_4348 : _GEN_4309; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4388 = _T_812 ? _GEN_4349 : _GEN_4310; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4389 = _T_812 ? _GEN_4350 : _GEN_4311; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4390 = _T_812 ? _GEN_4351 : _GEN_4312; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4391 = _T_812 ? _GEN_4352 : _GEN_4313; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4392 = _T_812 ? _GEN_4353 : _GEN_4314; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4393 = _T_812 ? _GEN_4354 : _GEN_4315; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4394 = _T_812 ? _GEN_4355 : _GEN_4316; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4395 = _T_812 ? _GEN_4356 : _GEN_4317; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4396 = _T_812 ? _GEN_4357 : _GEN_4318; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4397 = _T_812 ? _GEN_4358 : _GEN_4319; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4398 = _T_812 ? _GEN_4359 : _GEN_4320; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4399 = _T_812 ? _GEN_4360 : _GEN_4321; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4400 = _T_812 ? _GEN_4361 : _GEN_4322; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4401 = _T_812 ? _GEN_4362 : _GEN_4323; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_4402 = _T_812 ? _GEN_4363 : _GEN_4324; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [6:0] _funct7_T_11 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_56 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_824 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_50 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_128 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:65]
  wire [31:0] _now_reg_rs2_22 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_129 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:87]
  wire [63:0] _next_reg_T_130 = $signed(_T_300) * $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:72]
  wire [63:0] _next_reg_T_131 = $signed(_T_300) * $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:95]
  wire [31:0] _next_reg_T_132 = _next_reg_T_131[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:101]
  wire [31:0] _next_reg_rd_35 = _next_reg_T_131[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:101]
  wire [31:0] _GEN_4403 = 5'h0 == rd ? _next_reg_T_131[63:32] : _GEN_4371; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4404 = 5'h1 == rd ? _next_reg_T_131[63:32] : _GEN_4372; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4405 = 5'h2 == rd ? _next_reg_T_131[63:32] : _GEN_4373; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4406 = 5'h3 == rd ? _next_reg_T_131[63:32] : _GEN_4374; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4407 = 5'h4 == rd ? _next_reg_T_131[63:32] : _GEN_4375; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4408 = 5'h5 == rd ? _next_reg_T_131[63:32] : _GEN_4376; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4409 = 5'h6 == rd ? _next_reg_T_131[63:32] : _GEN_4377; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4410 = 5'h7 == rd ? _next_reg_T_131[63:32] : _GEN_4378; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4411 = 5'h8 == rd ? _next_reg_T_131[63:32] : _GEN_4379; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4412 = 5'h9 == rd ? _next_reg_T_131[63:32] : _GEN_4380; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4413 = 5'ha == rd ? _next_reg_T_131[63:32] : _GEN_4381; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4414 = 5'hb == rd ? _next_reg_T_131[63:32] : _GEN_4382; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4415 = 5'hc == rd ? _next_reg_T_131[63:32] : _GEN_4383; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4416 = 5'hd == rd ? _next_reg_T_131[63:32] : _GEN_4384; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4417 = 5'he == rd ? _next_reg_T_131[63:32] : _GEN_4385; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4418 = 5'hf == rd ? _next_reg_T_131[63:32] : _GEN_4386; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4419 = 5'h10 == rd ? _next_reg_T_131[63:32] : _GEN_4387; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4420 = 5'h11 == rd ? _next_reg_T_131[63:32] : _GEN_4388; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4421 = 5'h12 == rd ? _next_reg_T_131[63:32] : _GEN_4389; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4422 = 5'h13 == rd ? _next_reg_T_131[63:32] : _GEN_4390; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4423 = 5'h14 == rd ? _next_reg_T_131[63:32] : _GEN_4391; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4424 = 5'h15 == rd ? _next_reg_T_131[63:32] : _GEN_4392; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4425 = 5'h16 == rd ? _next_reg_T_131[63:32] : _GEN_4393; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4426 = 5'h17 == rd ? _next_reg_T_131[63:32] : _GEN_4394; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4427 = 5'h18 == rd ? _next_reg_T_131[63:32] : _GEN_4395; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4428 = 5'h19 == rd ? _next_reg_T_131[63:32] : _GEN_4396; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4429 = 5'h1a == rd ? _next_reg_T_131[63:32] : _GEN_4397; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4430 = 5'h1b == rd ? _next_reg_T_131[63:32] : _GEN_4398; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4431 = 5'h1c == rd ? _next_reg_T_131[63:32] : _GEN_4399; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4432 = 5'h1d == rd ? _next_reg_T_131[63:32] : _GEN_4400; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4433 = 5'h1e == rd ? _next_reg_T_131[63:32] : _GEN_4401; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_4434 = 5'h1f == rd ? _next_reg_T_131[63:32] : _GEN_4402; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [6:0] _GEN_4436 = _T_819 ? inst[31:25] : _GEN_4365; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4439 = _T_819 ? inst[14:12] : _GEN_4368; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4441 = _T_819 ? inst[6:0] : _GEN_4370; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4442 = _T_819 ? _GEN_4403 : _GEN_4371; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4443 = _T_819 ? _GEN_4404 : _GEN_4372; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4444 = _T_819 ? _GEN_4405 : _GEN_4373; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4445 = _T_819 ? _GEN_4406 : _GEN_4374; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4446 = _T_819 ? _GEN_4407 : _GEN_4375; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4447 = _T_819 ? _GEN_4408 : _GEN_4376; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4448 = _T_819 ? _GEN_4409 : _GEN_4377; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4449 = _T_819 ? _GEN_4410 : _GEN_4378; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4450 = _T_819 ? _GEN_4411 : _GEN_4379; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4451 = _T_819 ? _GEN_4412 : _GEN_4380; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4452 = _T_819 ? _GEN_4413 : _GEN_4381; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4453 = _T_819 ? _GEN_4414 : _GEN_4382; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4454 = _T_819 ? _GEN_4415 : _GEN_4383; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4455 = _T_819 ? _GEN_4416 : _GEN_4384; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4456 = _T_819 ? _GEN_4417 : _GEN_4385; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4457 = _T_819 ? _GEN_4418 : _GEN_4386; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4458 = _T_819 ? _GEN_4419 : _GEN_4387; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4459 = _T_819 ? _GEN_4420 : _GEN_4388; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4460 = _T_819 ? _GEN_4421 : _GEN_4389; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4461 = _T_819 ? _GEN_4422 : _GEN_4390; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4462 = _T_819 ? _GEN_4423 : _GEN_4391; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4463 = _T_819 ? _GEN_4424 : _GEN_4392; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4464 = _T_819 ? _GEN_4425 : _GEN_4393; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4465 = _T_819 ? _GEN_4426 : _GEN_4394; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4466 = _T_819 ? _GEN_4427 : _GEN_4395; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4467 = _T_819 ? _GEN_4428 : _GEN_4396; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4468 = _T_819 ? _GEN_4429 : _GEN_4397; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4469 = _T_819 ? _GEN_4430 : _GEN_4398; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4470 = _T_819 ? _GEN_4431 : _GEN_4399; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4471 = _T_819 ? _GEN_4432 : _GEN_4400; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4472 = _T_819 ? _GEN_4433 : _GEN_4401; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_4473 = _T_819 ? _GEN_4434 : _GEN_4402; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [6:0] _funct7_T_12 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_57 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_831 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_51 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_133 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:65]
  wire [31:0] _now_reg_rs2_23 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_134 = {1'b0,$signed(_GEN_840)}; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [64:0] _next_reg_T_135 = $signed(_T_300) * $signed(_next_reg_T_134); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [63:0] _next_reg_T_136 = _next_reg_T_135[63:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [63:0] _next_reg_T_137 = _next_reg_T_135[63:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [63:0] _next_reg_T_138 = _next_reg_T_135[63:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:88]
  wire [31:0] _next_reg_T_139 = _next_reg_T_138[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:94]
  wire [31:0] _next_reg_rd_36 = _next_reg_T_138[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:94]
  wire [31:0] _GEN_4474 = 5'h0 == rd ? _next_reg_T_138[63:32] : _GEN_4442; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4475 = 5'h1 == rd ? _next_reg_T_138[63:32] : _GEN_4443; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4476 = 5'h2 == rd ? _next_reg_T_138[63:32] : _GEN_4444; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4477 = 5'h3 == rd ? _next_reg_T_138[63:32] : _GEN_4445; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4478 = 5'h4 == rd ? _next_reg_T_138[63:32] : _GEN_4446; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4479 = 5'h5 == rd ? _next_reg_T_138[63:32] : _GEN_4447; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4480 = 5'h6 == rd ? _next_reg_T_138[63:32] : _GEN_4448; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4481 = 5'h7 == rd ? _next_reg_T_138[63:32] : _GEN_4449; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4482 = 5'h8 == rd ? _next_reg_T_138[63:32] : _GEN_4450; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4483 = 5'h9 == rd ? _next_reg_T_138[63:32] : _GEN_4451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4484 = 5'ha == rd ? _next_reg_T_138[63:32] : _GEN_4452; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4485 = 5'hb == rd ? _next_reg_T_138[63:32] : _GEN_4453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4486 = 5'hc == rd ? _next_reg_T_138[63:32] : _GEN_4454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4487 = 5'hd == rd ? _next_reg_T_138[63:32] : _GEN_4455; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4488 = 5'he == rd ? _next_reg_T_138[63:32] : _GEN_4456; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4489 = 5'hf == rd ? _next_reg_T_138[63:32] : _GEN_4457; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4490 = 5'h10 == rd ? _next_reg_T_138[63:32] : _GEN_4458; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4491 = 5'h11 == rd ? _next_reg_T_138[63:32] : _GEN_4459; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4492 = 5'h12 == rd ? _next_reg_T_138[63:32] : _GEN_4460; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4493 = 5'h13 == rd ? _next_reg_T_138[63:32] : _GEN_4461; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4494 = 5'h14 == rd ? _next_reg_T_138[63:32] : _GEN_4462; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4495 = 5'h15 == rd ? _next_reg_T_138[63:32] : _GEN_4463; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4496 = 5'h16 == rd ? _next_reg_T_138[63:32] : _GEN_4464; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4497 = 5'h17 == rd ? _next_reg_T_138[63:32] : _GEN_4465; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4498 = 5'h18 == rd ? _next_reg_T_138[63:32] : _GEN_4466; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4499 = 5'h19 == rd ? _next_reg_T_138[63:32] : _GEN_4467; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4500 = 5'h1a == rd ? _next_reg_T_138[63:32] : _GEN_4468; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4501 = 5'h1b == rd ? _next_reg_T_138[63:32] : _GEN_4469; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4502 = 5'h1c == rd ? _next_reg_T_138[63:32] : _GEN_4470; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4503 = 5'h1d == rd ? _next_reg_T_138[63:32] : _GEN_4471; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4504 = 5'h1e == rd ? _next_reg_T_138[63:32] : _GEN_4472; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_4505 = 5'h1f == rd ? _next_reg_T_138[63:32] : _GEN_4473; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [6:0] _GEN_4507 = _T_826 ? inst[31:25] : _GEN_4436; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4510 = _T_826 ? inst[14:12] : _GEN_4439; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4512 = _T_826 ? inst[6:0] : _GEN_4441; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4513 = _T_826 ? _GEN_4474 : _GEN_4442; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4514 = _T_826 ? _GEN_4475 : _GEN_4443; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4515 = _T_826 ? _GEN_4476 : _GEN_4444; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4516 = _T_826 ? _GEN_4477 : _GEN_4445; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4517 = _T_826 ? _GEN_4478 : _GEN_4446; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4518 = _T_826 ? _GEN_4479 : _GEN_4447; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4519 = _T_826 ? _GEN_4480 : _GEN_4448; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4520 = _T_826 ? _GEN_4481 : _GEN_4449; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4521 = _T_826 ? _GEN_4482 : _GEN_4450; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4522 = _T_826 ? _GEN_4483 : _GEN_4451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4523 = _T_826 ? _GEN_4484 : _GEN_4452; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4524 = _T_826 ? _GEN_4485 : _GEN_4453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4525 = _T_826 ? _GEN_4486 : _GEN_4454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4526 = _T_826 ? _GEN_4487 : _GEN_4455; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4527 = _T_826 ? _GEN_4488 : _GEN_4456; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4528 = _T_826 ? _GEN_4489 : _GEN_4457; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4529 = _T_826 ? _GEN_4490 : _GEN_4458; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4530 = _T_826 ? _GEN_4491 : _GEN_4459; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4531 = _T_826 ? _GEN_4492 : _GEN_4460; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4532 = _T_826 ? _GEN_4493 : _GEN_4461; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4533 = _T_826 ? _GEN_4494 : _GEN_4462; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4534 = _T_826 ? _GEN_4495 : _GEN_4463; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4535 = _T_826 ? _GEN_4496 : _GEN_4464; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4536 = _T_826 ? _GEN_4497 : _GEN_4465; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4537 = _T_826 ? _GEN_4498 : _GEN_4466; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4538 = _T_826 ? _GEN_4499 : _GEN_4467; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4539 = _T_826 ? _GEN_4500 : _GEN_4468; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4540 = _T_826 ? _GEN_4501 : _GEN_4469; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4541 = _T_826 ? _GEN_4502 : _GEN_4470; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4542 = _T_826 ? _GEN_4503 : _GEN_4471; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4543 = _T_826 ? _GEN_4504 : _GEN_4472; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_4544 = _T_826 ? _GEN_4505 : _GEN_4473; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [6:0] _funct7_T_13 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_58 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_838 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_52 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_24 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _next_reg_T_140 = _GEN_31 * _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:65]
  wire [31:0] _next_reg_T_141 = _next_reg_T_126[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:80]
  wire [31:0] _next_reg_rd_37 = _next_reg_T_126[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:80]
  wire [31:0] _GEN_4545 = 5'h0 == rd ? _next_reg_T_126[63:32] : _GEN_4513; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4546 = 5'h1 == rd ? _next_reg_T_126[63:32] : _GEN_4514; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4547 = 5'h2 == rd ? _next_reg_T_126[63:32] : _GEN_4515; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4548 = 5'h3 == rd ? _next_reg_T_126[63:32] : _GEN_4516; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4549 = 5'h4 == rd ? _next_reg_T_126[63:32] : _GEN_4517; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4550 = 5'h5 == rd ? _next_reg_T_126[63:32] : _GEN_4518; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4551 = 5'h6 == rd ? _next_reg_T_126[63:32] : _GEN_4519; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4552 = 5'h7 == rd ? _next_reg_T_126[63:32] : _GEN_4520; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4553 = 5'h8 == rd ? _next_reg_T_126[63:32] : _GEN_4521; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4554 = 5'h9 == rd ? _next_reg_T_126[63:32] : _GEN_4522; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4555 = 5'ha == rd ? _next_reg_T_126[63:32] : _GEN_4523; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4556 = 5'hb == rd ? _next_reg_T_126[63:32] : _GEN_4524; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4557 = 5'hc == rd ? _next_reg_T_126[63:32] : _GEN_4525; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4558 = 5'hd == rd ? _next_reg_T_126[63:32] : _GEN_4526; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4559 = 5'he == rd ? _next_reg_T_126[63:32] : _GEN_4527; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4560 = 5'hf == rd ? _next_reg_T_126[63:32] : _GEN_4528; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4561 = 5'h10 == rd ? _next_reg_T_126[63:32] : _GEN_4529; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4562 = 5'h11 == rd ? _next_reg_T_126[63:32] : _GEN_4530; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4563 = 5'h12 == rd ? _next_reg_T_126[63:32] : _GEN_4531; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4564 = 5'h13 == rd ? _next_reg_T_126[63:32] : _GEN_4532; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4565 = 5'h14 == rd ? _next_reg_T_126[63:32] : _GEN_4533; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4566 = 5'h15 == rd ? _next_reg_T_126[63:32] : _GEN_4534; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4567 = 5'h16 == rd ? _next_reg_T_126[63:32] : _GEN_4535; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4568 = 5'h17 == rd ? _next_reg_T_126[63:32] : _GEN_4536; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4569 = 5'h18 == rd ? _next_reg_T_126[63:32] : _GEN_4537; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4570 = 5'h19 == rd ? _next_reg_T_126[63:32] : _GEN_4538; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4571 = 5'h1a == rd ? _next_reg_T_126[63:32] : _GEN_4539; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4572 = 5'h1b == rd ? _next_reg_T_126[63:32] : _GEN_4540; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4573 = 5'h1c == rd ? _next_reg_T_126[63:32] : _GEN_4541; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4574 = 5'h1d == rd ? _next_reg_T_126[63:32] : _GEN_4542; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4575 = 5'h1e == rd ? _next_reg_T_126[63:32] : _GEN_4543; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_4576 = 5'h1f == rd ? _next_reg_T_126[63:32] : _GEN_4544; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [6:0] _GEN_4578 = _T_833 ? inst[31:25] : _GEN_4507; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4581 = _T_833 ? inst[14:12] : _GEN_4510; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4583 = _T_833 ? inst[6:0] : _GEN_4512; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4584 = _T_833 ? _GEN_4545 : _GEN_4513; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4585 = _T_833 ? _GEN_4546 : _GEN_4514; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4586 = _T_833 ? _GEN_4547 : _GEN_4515; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4587 = _T_833 ? _GEN_4548 : _GEN_4516; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4588 = _T_833 ? _GEN_4549 : _GEN_4517; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4589 = _T_833 ? _GEN_4550 : _GEN_4518; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4590 = _T_833 ? _GEN_4551 : _GEN_4519; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4591 = _T_833 ? _GEN_4552 : _GEN_4520; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4592 = _T_833 ? _GEN_4553 : _GEN_4521; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4593 = _T_833 ? _GEN_4554 : _GEN_4522; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4594 = _T_833 ? _GEN_4555 : _GEN_4523; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4595 = _T_833 ? _GEN_4556 : _GEN_4524; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4596 = _T_833 ? _GEN_4557 : _GEN_4525; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4597 = _T_833 ? _GEN_4558 : _GEN_4526; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4598 = _T_833 ? _GEN_4559 : _GEN_4527; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4599 = _T_833 ? _GEN_4560 : _GEN_4528; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4600 = _T_833 ? _GEN_4561 : _GEN_4529; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4601 = _T_833 ? _GEN_4562 : _GEN_4530; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4602 = _T_833 ? _GEN_4563 : _GEN_4531; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4603 = _T_833 ? _GEN_4564 : _GEN_4532; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4604 = _T_833 ? _GEN_4565 : _GEN_4533; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4605 = _T_833 ? _GEN_4566 : _GEN_4534; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4606 = _T_833 ? _GEN_4567 : _GEN_4535; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4607 = _T_833 ? _GEN_4568 : _GEN_4536; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4608 = _T_833 ? _GEN_4569 : _GEN_4537; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4609 = _T_833 ? _GEN_4570 : _GEN_4538; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4610 = _T_833 ? _GEN_4571 : _GEN_4539; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4611 = _T_833 ? _GEN_4572 : _GEN_4540; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4612 = _T_833 ? _GEN_4573 : _GEN_4541; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4613 = _T_833 ? _GEN_4574 : _GEN_4542; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4614 = _T_833 ? _GEN_4575 : _GEN_4543; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_4615 = _T_833 ? _GEN_4576 : _GEN_4544; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [6:0] _funct7_T_14 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_59 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_845 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_53 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_142 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:16]
  wire [31:0] _now_reg_rs2_25 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_143 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:34]
  wire [32:0] _next_reg_T_144 = $signed(_T_300) / $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:23]
  wire [31:0] _next_reg_T_145 = _next_reg_T_144[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:41]
  wire [31:0] _now_reg_rs2_26 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_146 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:19]
  wire [31:0] _next_reg_T_147 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:99]
  wire [31:0] _next_reg_T_148 = 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:45]
  wire [32:0] _next_reg_T_149 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire [31:0] _next_reg_T_150 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire [31:0] _now_reg_rs1_54 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _next_reg_T_151 = _GEN_31 == _next_reg_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:18]
  wire [31:0] _next_reg_T_152 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:78]
  wire [31:0] _now_reg_rs2_27 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_153 = _GEN_840 == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:64]
  wire  _next_reg_T_154 = _GEN_31 == _next_reg_T_150 & _GEN_840 == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:52]
  wire [31:0] _next_reg_T_155 = 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:112]
  wire [32:0] _next_reg_T_156 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:89]
  wire [31:0] _next_reg_T_157 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:89]
  wire [31:0] _next_reg_T_158 = _next_reg_T_154 ? _next_reg_T_150 : _next_reg_T_144[31:0]; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_T_159 = _next_reg_T_146 ? 32'hffffffff : _next_reg_T_158; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_38 = _next_reg_T_146 ? 32'hffffffff : _next_reg_T_158; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_4616 = 5'h0 == rd ? _next_reg_T_159 : _GEN_4584; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4617 = 5'h1 == rd ? _next_reg_T_159 : _GEN_4585; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4618 = 5'h2 == rd ? _next_reg_T_159 : _GEN_4586; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4619 = 5'h3 == rd ? _next_reg_T_159 : _GEN_4587; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4620 = 5'h4 == rd ? _next_reg_T_159 : _GEN_4588; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4621 = 5'h5 == rd ? _next_reg_T_159 : _GEN_4589; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4622 = 5'h6 == rd ? _next_reg_T_159 : _GEN_4590; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4623 = 5'h7 == rd ? _next_reg_T_159 : _GEN_4591; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4624 = 5'h8 == rd ? _next_reg_T_159 : _GEN_4592; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4625 = 5'h9 == rd ? _next_reg_T_159 : _GEN_4593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4626 = 5'ha == rd ? _next_reg_T_159 : _GEN_4594; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4627 = 5'hb == rd ? _next_reg_T_159 : _GEN_4595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4628 = 5'hc == rd ? _next_reg_T_159 : _GEN_4596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4629 = 5'hd == rd ? _next_reg_T_159 : _GEN_4597; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4630 = 5'he == rd ? _next_reg_T_159 : _GEN_4598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4631 = 5'hf == rd ? _next_reg_T_159 : _GEN_4599; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4632 = 5'h10 == rd ? _next_reg_T_159 : _GEN_4600; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4633 = 5'h11 == rd ? _next_reg_T_159 : _GEN_4601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4634 = 5'h12 == rd ? _next_reg_T_159 : _GEN_4602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4635 = 5'h13 == rd ? _next_reg_T_159 : _GEN_4603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4636 = 5'h14 == rd ? _next_reg_T_159 : _GEN_4604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4637 = 5'h15 == rd ? _next_reg_T_159 : _GEN_4605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4638 = 5'h16 == rd ? _next_reg_T_159 : _GEN_4606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4639 = 5'h17 == rd ? _next_reg_T_159 : _GEN_4607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4640 = 5'h18 == rd ? _next_reg_T_159 : _GEN_4608; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4641 = 5'h19 == rd ? _next_reg_T_159 : _GEN_4609; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4642 = 5'h1a == rd ? _next_reg_T_159 : _GEN_4610; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4643 = 5'h1b == rd ? _next_reg_T_159 : _GEN_4611; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4644 = 5'h1c == rd ? _next_reg_T_159 : _GEN_4612; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4645 = 5'h1d == rd ? _next_reg_T_159 : _GEN_4613; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4646 = 5'h1e == rd ? _next_reg_T_159 : _GEN_4614; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_4647 = 5'h1f == rd ? _next_reg_T_159 : _GEN_4615; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [6:0] _GEN_4649 = _T_840 ? inst[31:25] : _GEN_4578; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4652 = _T_840 ? inst[14:12] : _GEN_4581; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4654 = _T_840 ? inst[6:0] : _GEN_4583; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4655 = _T_840 ? _GEN_4616 : _GEN_4584; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4656 = _T_840 ? _GEN_4617 : _GEN_4585; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4657 = _T_840 ? _GEN_4618 : _GEN_4586; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4658 = _T_840 ? _GEN_4619 : _GEN_4587; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4659 = _T_840 ? _GEN_4620 : _GEN_4588; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4660 = _T_840 ? _GEN_4621 : _GEN_4589; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4661 = _T_840 ? _GEN_4622 : _GEN_4590; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4662 = _T_840 ? _GEN_4623 : _GEN_4591; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4663 = _T_840 ? _GEN_4624 : _GEN_4592; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4664 = _T_840 ? _GEN_4625 : _GEN_4593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4665 = _T_840 ? _GEN_4626 : _GEN_4594; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4666 = _T_840 ? _GEN_4627 : _GEN_4595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4667 = _T_840 ? _GEN_4628 : _GEN_4596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4668 = _T_840 ? _GEN_4629 : _GEN_4597; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4669 = _T_840 ? _GEN_4630 : _GEN_4598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4670 = _T_840 ? _GEN_4631 : _GEN_4599; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4671 = _T_840 ? _GEN_4632 : _GEN_4600; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4672 = _T_840 ? _GEN_4633 : _GEN_4601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4673 = _T_840 ? _GEN_4634 : _GEN_4602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4674 = _T_840 ? _GEN_4635 : _GEN_4603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4675 = _T_840 ? _GEN_4636 : _GEN_4604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4676 = _T_840 ? _GEN_4637 : _GEN_4605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4677 = _T_840 ? _GEN_4638 : _GEN_4606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4678 = _T_840 ? _GEN_4639 : _GEN_4607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4679 = _T_840 ? _GEN_4640 : _GEN_4608; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4680 = _T_840 ? _GEN_4641 : _GEN_4609; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4681 = _T_840 ? _GEN_4642 : _GEN_4610; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4682 = _T_840 ? _GEN_4643 : _GEN_4611; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4683 = _T_840 ? _GEN_4644 : _GEN_4612; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4684 = _T_840 ? _GEN_4645 : _GEN_4613; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4685 = _T_840 ? _GEN_4646 : _GEN_4614; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_4686 = _T_840 ? _GEN_4647 : _GEN_4615; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [6:0] _funct7_T_15 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_60 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_852 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_55 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_28 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_160 = _GEN_31 / _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 58:15]
  wire [31:0] _now_reg_rs2_29 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_161 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 60:19]
  wire [31:0] _next_reg_T_162 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 60:40]
  wire [31:0] _next_reg_T_163 = _next_reg_T_146 ? 32'hffffffff : _next_reg_T_160; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_39 = _next_reg_T_146 ? 32'hffffffff : _next_reg_T_160; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_4687 = 5'h0 == rd ? _next_reg_T_163 : _GEN_4655; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4688 = 5'h1 == rd ? _next_reg_T_163 : _GEN_4656; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4689 = 5'h2 == rd ? _next_reg_T_163 : _GEN_4657; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4690 = 5'h3 == rd ? _next_reg_T_163 : _GEN_4658; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4691 = 5'h4 == rd ? _next_reg_T_163 : _GEN_4659; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4692 = 5'h5 == rd ? _next_reg_T_163 : _GEN_4660; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4693 = 5'h6 == rd ? _next_reg_T_163 : _GEN_4661; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4694 = 5'h7 == rd ? _next_reg_T_163 : _GEN_4662; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4695 = 5'h8 == rd ? _next_reg_T_163 : _GEN_4663; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4696 = 5'h9 == rd ? _next_reg_T_163 : _GEN_4664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4697 = 5'ha == rd ? _next_reg_T_163 : _GEN_4665; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4698 = 5'hb == rd ? _next_reg_T_163 : _GEN_4666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4699 = 5'hc == rd ? _next_reg_T_163 : _GEN_4667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4700 = 5'hd == rd ? _next_reg_T_163 : _GEN_4668; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4701 = 5'he == rd ? _next_reg_T_163 : _GEN_4669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4702 = 5'hf == rd ? _next_reg_T_163 : _GEN_4670; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4703 = 5'h10 == rd ? _next_reg_T_163 : _GEN_4671; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4704 = 5'h11 == rd ? _next_reg_T_163 : _GEN_4672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4705 = 5'h12 == rd ? _next_reg_T_163 : _GEN_4673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4706 = 5'h13 == rd ? _next_reg_T_163 : _GEN_4674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4707 = 5'h14 == rd ? _next_reg_T_163 : _GEN_4675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4708 = 5'h15 == rd ? _next_reg_T_163 : _GEN_4676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4709 = 5'h16 == rd ? _next_reg_T_163 : _GEN_4677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4710 = 5'h17 == rd ? _next_reg_T_163 : _GEN_4678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4711 = 5'h18 == rd ? _next_reg_T_163 : _GEN_4679; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4712 = 5'h19 == rd ? _next_reg_T_163 : _GEN_4680; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4713 = 5'h1a == rd ? _next_reg_T_163 : _GEN_4681; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4714 = 5'h1b == rd ? _next_reg_T_163 : _GEN_4682; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4715 = 5'h1c == rd ? _next_reg_T_163 : _GEN_4683; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4716 = 5'h1d == rd ? _next_reg_T_163 : _GEN_4684; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4717 = 5'h1e == rd ? _next_reg_T_163 : _GEN_4685; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_4718 = 5'h1f == rd ? _next_reg_T_163 : _GEN_4686; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [6:0] _GEN_4720 = _T_847 ? inst[31:25] : _GEN_4649; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4723 = _T_847 ? inst[14:12] : _GEN_4652; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4725 = _T_847 ? inst[6:0] : _GEN_4654; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4726 = _T_847 ? _GEN_4687 : _GEN_4655; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4727 = _T_847 ? _GEN_4688 : _GEN_4656; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4728 = _T_847 ? _GEN_4689 : _GEN_4657; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4729 = _T_847 ? _GEN_4690 : _GEN_4658; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4730 = _T_847 ? _GEN_4691 : _GEN_4659; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4731 = _T_847 ? _GEN_4692 : _GEN_4660; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4732 = _T_847 ? _GEN_4693 : _GEN_4661; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4733 = _T_847 ? _GEN_4694 : _GEN_4662; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4734 = _T_847 ? _GEN_4695 : _GEN_4663; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4735 = _T_847 ? _GEN_4696 : _GEN_4664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4736 = _T_847 ? _GEN_4697 : _GEN_4665; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4737 = _T_847 ? _GEN_4698 : _GEN_4666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4738 = _T_847 ? _GEN_4699 : _GEN_4667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4739 = _T_847 ? _GEN_4700 : _GEN_4668; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4740 = _T_847 ? _GEN_4701 : _GEN_4669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4741 = _T_847 ? _GEN_4702 : _GEN_4670; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4742 = _T_847 ? _GEN_4703 : _GEN_4671; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4743 = _T_847 ? _GEN_4704 : _GEN_4672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4744 = _T_847 ? _GEN_4705 : _GEN_4673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4745 = _T_847 ? _GEN_4706 : _GEN_4674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4746 = _T_847 ? _GEN_4707 : _GEN_4675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4747 = _T_847 ? _GEN_4708 : _GEN_4676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4748 = _T_847 ? _GEN_4709 : _GEN_4677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4749 = _T_847 ? _GEN_4710 : _GEN_4678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4750 = _T_847 ? _GEN_4711 : _GEN_4679; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4751 = _T_847 ? _GEN_4712 : _GEN_4680; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4752 = _T_847 ? _GEN_4713 : _GEN_4681; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4753 = _T_847 ? _GEN_4714 : _GEN_4682; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4754 = _T_847 ? _GEN_4715 : _GEN_4683; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4755 = _T_847 ? _GEN_4716 : _GEN_4684; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4756 = _T_847 ? _GEN_4717 : _GEN_4685; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_4757 = _T_847 ? _GEN_4718 : _GEN_4686; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [6:0] _funct7_T_16 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_61 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_859 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_56 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_164 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:16]
  wire [31:0] _now_reg_rs2_30 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_165 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:34]
  wire [31:0] _next_reg_T_166 = $signed(_T_300) % $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:23]
  wire [31:0] _next_reg_T_167 = $signed(_T_300) % $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:42]
  wire [31:0] _now_reg_rs2_31 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_168 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 68:19]
  wire [31:0] _next_reg_T_169 = 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:45]
  wire [32:0] _next_reg_T_170 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:22]
  wire [31:0] _next_reg_T_171 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:22]
  wire [31:0] _now_reg_rs1_57 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _next_reg_T_172 = _GEN_31 == _next_reg_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:18]
  wire [31:0] _next_reg_T_173 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:78]
  wire [31:0] _now_reg_rs2_32 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_174 = _GEN_840 == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:64]
  wire  _next_reg_T_175 = _next_reg_T_151 & _next_reg_T_153; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:52]
  wire [31:0] _next_reg_T_176 = _next_reg_T_154 ? 32'h0 : _next_reg_T_167; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _now_reg_rs1_58 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_177 = _next_reg_T_146 ? _GEN_31 : _next_reg_T_176; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_40 = _next_reg_T_146 ? _GEN_31 : _next_reg_T_176; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_4758 = 5'h0 == rd ? _next_reg_T_177 : _GEN_4726; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4759 = 5'h1 == rd ? _next_reg_T_177 : _GEN_4727; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4760 = 5'h2 == rd ? _next_reg_T_177 : _GEN_4728; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4761 = 5'h3 == rd ? _next_reg_T_177 : _GEN_4729; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4762 = 5'h4 == rd ? _next_reg_T_177 : _GEN_4730; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4763 = 5'h5 == rd ? _next_reg_T_177 : _GEN_4731; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4764 = 5'h6 == rd ? _next_reg_T_177 : _GEN_4732; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4765 = 5'h7 == rd ? _next_reg_T_177 : _GEN_4733; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4766 = 5'h8 == rd ? _next_reg_T_177 : _GEN_4734; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4767 = 5'h9 == rd ? _next_reg_T_177 : _GEN_4735; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4768 = 5'ha == rd ? _next_reg_T_177 : _GEN_4736; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4769 = 5'hb == rd ? _next_reg_T_177 : _GEN_4737; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4770 = 5'hc == rd ? _next_reg_T_177 : _GEN_4738; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4771 = 5'hd == rd ? _next_reg_T_177 : _GEN_4739; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4772 = 5'he == rd ? _next_reg_T_177 : _GEN_4740; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4773 = 5'hf == rd ? _next_reg_T_177 : _GEN_4741; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4774 = 5'h10 == rd ? _next_reg_T_177 : _GEN_4742; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4775 = 5'h11 == rd ? _next_reg_T_177 : _GEN_4743; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4776 = 5'h12 == rd ? _next_reg_T_177 : _GEN_4744; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4777 = 5'h13 == rd ? _next_reg_T_177 : _GEN_4745; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4778 = 5'h14 == rd ? _next_reg_T_177 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4779 = 5'h15 == rd ? _next_reg_T_177 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4780 = 5'h16 == rd ? _next_reg_T_177 : _GEN_4748; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4781 = 5'h17 == rd ? _next_reg_T_177 : _GEN_4749; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4782 = 5'h18 == rd ? _next_reg_T_177 : _GEN_4750; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4783 = 5'h19 == rd ? _next_reg_T_177 : _GEN_4751; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4784 = 5'h1a == rd ? _next_reg_T_177 : _GEN_4752; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4785 = 5'h1b == rd ? _next_reg_T_177 : _GEN_4753; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4786 = 5'h1c == rd ? _next_reg_T_177 : _GEN_4754; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4787 = 5'h1d == rd ? _next_reg_T_177 : _GEN_4755; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4788 = 5'h1e == rd ? _next_reg_T_177 : _GEN_4756; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_4789 = 5'h1f == rd ? _next_reg_T_177 : _GEN_4757; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [6:0] _GEN_4791 = _T_854 ? inst[31:25] : _GEN_4720; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4794 = _T_854 ? inst[14:12] : _GEN_4723; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4796 = _T_854 ? inst[6:0] : _GEN_4725; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4797 = _T_854 ? _GEN_4758 : _GEN_4726; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4798 = _T_854 ? _GEN_4759 : _GEN_4727; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4799 = _T_854 ? _GEN_4760 : _GEN_4728; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4800 = _T_854 ? _GEN_4761 : _GEN_4729; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4801 = _T_854 ? _GEN_4762 : _GEN_4730; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4802 = _T_854 ? _GEN_4763 : _GEN_4731; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4803 = _T_854 ? _GEN_4764 : _GEN_4732; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4804 = _T_854 ? _GEN_4765 : _GEN_4733; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4805 = _T_854 ? _GEN_4766 : _GEN_4734; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4806 = _T_854 ? _GEN_4767 : _GEN_4735; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4807 = _T_854 ? _GEN_4768 : _GEN_4736; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4808 = _T_854 ? _GEN_4769 : _GEN_4737; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4809 = _T_854 ? _GEN_4770 : _GEN_4738; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4810 = _T_854 ? _GEN_4771 : _GEN_4739; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4811 = _T_854 ? _GEN_4772 : _GEN_4740; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4812 = _T_854 ? _GEN_4773 : _GEN_4741; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4813 = _T_854 ? _GEN_4774 : _GEN_4742; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4814 = _T_854 ? _GEN_4775 : _GEN_4743; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4815 = _T_854 ? _GEN_4776 : _GEN_4744; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4816 = _T_854 ? _GEN_4777 : _GEN_4745; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4817 = _T_854 ? _GEN_4778 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4818 = _T_854 ? _GEN_4779 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4819 = _T_854 ? _GEN_4780 : _GEN_4748; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4820 = _T_854 ? _GEN_4781 : _GEN_4749; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4821 = _T_854 ? _GEN_4782 : _GEN_4750; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4822 = _T_854 ? _GEN_4783 : _GEN_4751; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4823 = _T_854 ? _GEN_4784 : _GEN_4752; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4824 = _T_854 ? _GEN_4785 : _GEN_4753; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4825 = _T_854 ? _GEN_4786 : _GEN_4754; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4826 = _T_854 ? _GEN_4787 : _GEN_4755; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4827 = _T_854 ? _GEN_4788 : _GEN_4756; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_4828 = _T_854 ? _GEN_4789 : _GEN_4757; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [6:0] _funct7_T_17 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_62 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_866 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_59 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_33 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_178 = _GEN_31 % _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 75:15]
  wire [31:0] _now_reg_rs2_34 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_179 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 77:19]
  wire [31:0] _now_reg_rs1_60 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_180 = _next_reg_T_146 ? _GEN_31 : _next_reg_T_178; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_41 = _next_reg_T_146 ? _GEN_31 : _next_reg_T_178; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_4829 = 5'h0 == rd ? _next_reg_T_180 : _GEN_4797; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4830 = 5'h1 == rd ? _next_reg_T_180 : _GEN_4798; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4831 = 5'h2 == rd ? _next_reg_T_180 : _GEN_4799; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4832 = 5'h3 == rd ? _next_reg_T_180 : _GEN_4800; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4833 = 5'h4 == rd ? _next_reg_T_180 : _GEN_4801; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4834 = 5'h5 == rd ? _next_reg_T_180 : _GEN_4802; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4835 = 5'h6 == rd ? _next_reg_T_180 : _GEN_4803; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4836 = 5'h7 == rd ? _next_reg_T_180 : _GEN_4804; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4837 = 5'h8 == rd ? _next_reg_T_180 : _GEN_4805; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4838 = 5'h9 == rd ? _next_reg_T_180 : _GEN_4806; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4839 = 5'ha == rd ? _next_reg_T_180 : _GEN_4807; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4840 = 5'hb == rd ? _next_reg_T_180 : _GEN_4808; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4841 = 5'hc == rd ? _next_reg_T_180 : _GEN_4809; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4842 = 5'hd == rd ? _next_reg_T_180 : _GEN_4810; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4843 = 5'he == rd ? _next_reg_T_180 : _GEN_4811; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4844 = 5'hf == rd ? _next_reg_T_180 : _GEN_4812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4845 = 5'h10 == rd ? _next_reg_T_180 : _GEN_4813; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4846 = 5'h11 == rd ? _next_reg_T_180 : _GEN_4814; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4847 = 5'h12 == rd ? _next_reg_T_180 : _GEN_4815; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4848 = 5'h13 == rd ? _next_reg_T_180 : _GEN_4816; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4849 = 5'h14 == rd ? _next_reg_T_180 : _GEN_4817; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4850 = 5'h15 == rd ? _next_reg_T_180 : _GEN_4818; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4851 = 5'h16 == rd ? _next_reg_T_180 : _GEN_4819; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4852 = 5'h17 == rd ? _next_reg_T_180 : _GEN_4820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4853 = 5'h18 == rd ? _next_reg_T_180 : _GEN_4821; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4854 = 5'h19 == rd ? _next_reg_T_180 : _GEN_4822; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4855 = 5'h1a == rd ? _next_reg_T_180 : _GEN_4823; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4856 = 5'h1b == rd ? _next_reg_T_180 : _GEN_4824; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4857 = 5'h1c == rd ? _next_reg_T_180 : _GEN_4825; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4858 = 5'h1d == rd ? _next_reg_T_180 : _GEN_4826; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4859 = 5'h1e == rd ? _next_reg_T_180 : _GEN_4827; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_4860 = 5'h1f == rd ? _next_reg_T_180 : _GEN_4828; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [6:0] _GEN_4862 = _T_861 ? inst[31:25] : _GEN_4791; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4865 = _T_861 ? inst[14:12] : _GEN_4794; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4867 = _T_861 ? inst[6:0] : _GEN_4796; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_4868 = _T_861 ? _GEN_4829 : _GEN_4797; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4869 = _T_861 ? _GEN_4830 : _GEN_4798; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4870 = _T_861 ? _GEN_4831 : _GEN_4799; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4871 = _T_861 ? _GEN_4832 : _GEN_4800; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4872 = _T_861 ? _GEN_4833 : _GEN_4801; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4873 = _T_861 ? _GEN_4834 : _GEN_4802; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4874 = _T_861 ? _GEN_4835 : _GEN_4803; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4875 = _T_861 ? _GEN_4836 : _GEN_4804; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4876 = _T_861 ? _GEN_4837 : _GEN_4805; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4877 = _T_861 ? _GEN_4838 : _GEN_4806; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4878 = _T_861 ? _GEN_4839 : _GEN_4807; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4879 = _T_861 ? _GEN_4840 : _GEN_4808; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4880 = _T_861 ? _GEN_4841 : _GEN_4809; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4881 = _T_861 ? _GEN_4842 : _GEN_4810; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4882 = _T_861 ? _GEN_4843 : _GEN_4811; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4883 = _T_861 ? _GEN_4844 : _GEN_4812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4884 = _T_861 ? _GEN_4845 : _GEN_4813; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4885 = _T_861 ? _GEN_4846 : _GEN_4814; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4886 = _T_861 ? _GEN_4847 : _GEN_4815; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4887 = _T_861 ? _GEN_4848 : _GEN_4816; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4888 = _T_861 ? _GEN_4849 : _GEN_4817; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4889 = _T_861 ? _GEN_4850 : _GEN_4818; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4890 = _T_861 ? _GEN_4851 : _GEN_4819; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4891 = _T_861 ? _GEN_4852 : _GEN_4820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4892 = _T_861 ? _GEN_4853 : _GEN_4821; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4893 = _T_861 ? _GEN_4854 : _GEN_4822; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4894 = _T_861 ? _GEN_4855 : _GEN_4823; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4895 = _T_861 ? _GEN_4856 : _GEN_4824; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4896 = _T_861 ? _GEN_4857 : _GEN_4825; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4897 = _T_861 ? _GEN_4858 : _GEN_4826; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4898 = _T_861 ? _GEN_4859 : _GEN_4827; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_4899 = _T_861 ? _GEN_4860 : _GEN_4828; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [2:0] _funct3_T_63 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_872 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  mstatusOld_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [7:0] mstatusOld_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [31:0] _mstatusNew_WIRE_1 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusNew_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_1 = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_5 = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_8 = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_13 = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [7:0] mstatusNew_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusOld_WIRE_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_8 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _next_internal_privilegeMode_T = {1'h0,mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 125:41]
  wire  _mstatusNew_WIRE_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusOld_WIRE_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_5 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusNew_sie = illegalSret | illegalSModeSret ? mstatusOld_sie : mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 124:35]
  wire  _GEN_4902 = mstatusNew_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 124:35]
  wire  _mstatusNew_WIRE_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] next_csr_mstatus_lo_lo_lo = {mstatusNew_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_4 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_3 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi = {mstatusOld_pad2,mstatusOld_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_2 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [2:0] next_csr_mstatus_lo_lo_hi = {mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [4:0] next_csr_mstatus_lo_lo = {mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3,mstatusNew_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_6 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_spie = illegalSret | illegalSModeSret ? mstatusOld_spie : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 126:35]
  wire  _GEN_4904 = mstatusNew_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 126:35]
  wire [1:0] next_csr_mstatus_lo_hi_lo = {mstatusOld_ube,mstatusNew_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [1:0] _mstatusNew_WIRE_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_9 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_spp = (illegalSret | illegalSModeSret) & mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 127:35]
  wire  _GEN_4905 = mstatusNew_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 127:35]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi = {mstatusOld_vs,mstatusNew_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_7 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [3:0] next_csr_mstatus_lo_hi_hi = {mstatusOld_vs,mstatusNew_spp,mstatusOld_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [5:0] next_csr_mstatus_lo_hi = {mstatusOld_vs,mstatusNew_spp,mstatusOld_mpie,mstatusOld_ube,mstatusNew_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [10:0] next_csr_mstatus_lo = {mstatusOld_vs,mstatusNew_spp,mstatusOld_mpie,mstatusOld_ube,mstatusNew_spie,
    mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3,mstatusNew_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [1:0] _mstatusNew_WIRE_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_11 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_WIRE_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_10 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [3:0] next_csr_mstatus_hi_lo_lo = {mstatusOld_fs,mstatusOld_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_14 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mprv = (illegalSret | illegalSModeSret) & mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 128:35]
  wire  _GEN_4906 = mstatusNew_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 128:35]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi = {mstatusOld_sum,mstatusNew_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [1:0] _mstatusNew_WIRE_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_12 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [3:0] next_csr_mstatus_hi_lo_hi = {mstatusOld_sum,mstatusNew_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [7:0] next_csr_mstatus_hi_lo = {mstatusOld_sum,mstatusNew_mprv,mstatusOld_xs,mstatusOld_fs,mstatusOld_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_17 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_16 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_15 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [2:0] next_csr_mstatus_hi_hi_lo = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_20 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [7:0] _mstatusNew_WIRE_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [7:0] _mstatusNew_T_19 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_18 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [9:0] next_csr_mstatus_hi_hi_hi = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [12:0] next_csr_mstatus_hi_hi = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [20:0] next_csr_mstatus_hi = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [31:0] _next_csr_mstatus_T = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo,next_csr_mstatus_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _GEN_4901 = illegalSret | illegalSModeSret | _GEN_2540; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_4919 = _T_868 ? _GEN_4901 : _GEN_2540; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire  _GEN_4931 = io_now_internal_privilegeMode == 2'h3 ? _GEN_4919 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_4945 = _T_875 ? _GEN_4931 : _GEN_4919; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_4961 = isIllegalAccess_5 | ~has_15 | _GEN_4945; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5051 = has_15 ? _GEN_4961 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5095 = _T_1089 ? _GEN_5051 : _GEN_4961; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire  _GEN_5105 = _T_894 ? _GEN_5095 : _GEN_4945; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire  _GEN_5149 = isIllegalAccess_4 | ~has_15 | _GEN_5105; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5211 = has_15 ? _GEN_5149 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5223 = _T_1090 ? _GEN_5211 : _GEN_5149; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire  _GEN_5267 = _T_1049 ? _GEN_5223 : _GEN_5149; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire  _GEN_5277 = _T_927 ? _GEN_5267 : _GEN_5105; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire  _GEN_5321 = isIllegalAccess_5 | ~has_15 | _GEN_5277; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5383 = has_15 ? _GEN_5321 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5395 = _T_1090 ? _GEN_5383 : _GEN_5321; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire  _GEN_5439 = _T_1089 ? _GEN_5395 : _GEN_5321; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire  _GEN_5449 = _T_967 ? _GEN_5439 : _GEN_5277; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire  _GEN_5493 = isIllegalAccess_5 | ~has_15 | _GEN_5449; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5583 = has_15 ? _GEN_5493 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5627 = _T_1089 ? _GEN_5583 : _GEN_5493; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire  _GEN_5637 = _T_1007 ? _GEN_5627 : _GEN_5449; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire  _GEN_5681 = isIllegalAccess_4 | ~has_15 | _GEN_5637; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5743 = has_15 ? _GEN_5681 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5755 = _T_1090 ? _GEN_5743 : _GEN_5681; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire  _GEN_5799 = ~isIllegalWrite_4 ? _GEN_5755 : _GEN_5681; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire  _GEN_5809 = _T_1041 ? _GEN_5799 : _GEN_5637; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire  _GEN_5853 = isIllegalAccess_5 | ~has_15 | _GEN_5809; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5915 = has_15 ? _GEN_5853 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5927 = rs1 != 5'h0 ? _GEN_5915 : _GEN_5853; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire  _GEN_5971 = ~isIllegalWrite_5 ? _GEN_5927 : _GEN_5853; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire  _GEN_5981 = _T_1082 ? _GEN_5971 : _GEN_5809; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire  _GEN_6026 = illegalInstruction | _GEN_5981; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 145:33]
  wire  raiseExceptionIntr = io_valid & _GEN_6026; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire  _GEN_6154 = raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [31:0] now_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _delegS_T = io_now_csr_medeleg >> exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:24]
  wire  _delegS_T_1 = _delegS_T[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:24]
  wire  _delegS_T_2 = io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:70]
  wire  delegS = _delegS_T[0] & io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:39]
  wire [7:0] now_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_1123 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] now_csr_sepc = io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6041 = 8'h20 == io_now_csr_MXLEN ? io_now_pc : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 254:35]
  wire [31:0] _GEN_6076 = delegS ? _GEN_6041 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_6093 = raiseExceptionIntr ? _GEN_6076 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_sepc = io_valid ? _GEN_6093 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6205 = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _retTarget_T = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [1:0] _GEN_4903 = illegalSret | illegalSModeSret ? io_now_internal_privilegeMode : _next_internal_privilegeMode_T
    ; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 125:35]
  wire [31:0] _GEN_4907 = illegalSret | illegalSModeSret ? io_now_csr_mstatus : _next_csr_mstatus_T; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 129:35]
  wire [31:0] _GEN_4908 = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  _GEN_4909 = illegalSret | illegalSModeSret ? _GEN_2936 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 132:25]
  wire [31:0] _GEN_4910 = illegalSret | illegalSModeSret ? _GEN_2937 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 133:25]
  wire [2:0] _GEN_4914 = _T_868 ? inst[14:12] : _GEN_4865; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4916 = _T_868 ? inst[6:0] : _GEN_4867; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [1:0] _GEN_4920 = _T_868 ? _GEN_4903 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_4921 = _T_868 ? _GEN_4907 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_4922 = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  _GEN_4923 = _T_868 ? _GEN_4909 : _GEN_2936; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_4924 = _T_868 ? _GEN_4910 : _GEN_2937; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [2:0] _funct3_T_64 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_879 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _mstatusOld_WIRE_3 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusOld_1_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [7:0] mstatusOld_1_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [31:0] _mstatusNew_WIRE_3 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusNew_1_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_24 = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_28 = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_31 = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [7:0] mstatusNew_1_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_22 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_21 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_lo_lo_lo_1 = {mstatusOld_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_25 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusOld_WIRE_2_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_28 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusNew_1_mie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_1 = {mstatusOld_pad2,mstatusOld_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_23 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [2:0] next_csr_mstatus_lo_lo_hi_1 = {mstatusOld_pad2,mstatusOld_mpie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [4:0] next_csr_mstatus_lo_lo_1 = {mstatusOld_pad2,mstatusOld_mpie,mstatusOld_pad3,mstatusOld_sie,mstatusOld_pad4}
    ; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_27 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_26 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_lo_hi_lo_1 = {mstatusOld_ube,mstatusOld_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [1:0] _mstatusNew_WIRE_2_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_30 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_29 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_1 = {mstatusOld_vs,mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  mstatusNew_1_mpie = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:32 93:35]
  wire [3:0] next_csr_mstatus_lo_hi_hi_1 = {mstatusOld_vs,mstatusOld_spp,1'h1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [5:0] next_csr_mstatus_lo_hi_1 = {mstatusOld_vs,mstatusOld_spp,1'h1,mstatusOld_ube,mstatusOld_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [10:0] next_csr_mstatus_lo_1 = {mstatusOld_vs,mstatusOld_spp,1'h1,mstatusOld_ube,mstatusOld_spie,mstatusOld_pad2,
    mstatusOld_mpie,mstatusOld_pad3,mstatusOld_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [1:0] _mstatusNew_WIRE_2_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_32 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_mpp = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:32 96:24]
  wire [3:0] next_csr_mstatus_hi_lo_lo_1 = {mstatusOld_fs,2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_35 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_34 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_1 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [1:0] _mstatusNew_WIRE_2_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_33 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [3:0] next_csr_mstatus_hi_lo_hi_1 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [7:0] next_csr_mstatus_hi_lo_1 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_38 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_37 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_1 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_36 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [2:0] next_csr_mstatus_hi_hi_lo_1 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_41 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [7:0] _mstatusNew_WIRE_2_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [7:0] _mstatusNew_T_40 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_1 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_39 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [9:0] next_csr_mstatus_hi_hi_hi_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [12:0] next_csr_mstatus_hi_hi_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [20:0] next_csr_mstatus_hi_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [31:0] _next_csr_mstatus_T_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_1,next_csr_mstatus_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _T_1116 = csrAddr == 12'h341; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] now_csr_mepc = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _next_csr_mepc_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mepc_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire  _T_1091 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_1092 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [7:0] now_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_1093 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _rData_T_20 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _rData_T_21 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _rData_T_22 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _rData_T_23 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire  _has_T_404 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_402 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_400 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_398 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_396 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_394 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_392 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_390 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_388 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_386 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_384 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_382 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_380 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_378 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_379 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_381 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_383 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_385 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_387 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_389 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_391 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_393 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_395 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_397 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_399 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_401 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_403 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  has_14 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _nowCSR_T_107 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_105 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mcause = io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_103 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_101 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mie = io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_99 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mip = io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_97 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mcounteren = io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_95 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mtvec = io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_93 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mscratch = io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_91 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_89 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_87 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_85 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_83 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] now_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _nowCSR_T_81 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_82 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_84 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_86 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_88 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_90 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_92 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_94 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_96 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_98 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_100 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_102 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_104 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_106 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] nowCSR_3 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _rData_T_18 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _rmask_T_163 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_136 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_161 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_135 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_159 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_134 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_157 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_133 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_155 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_132 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_153 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_131 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_151 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_130 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_149 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_129 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_147 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_128 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_145 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_127 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_143 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_126 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_141 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_125 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_139 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_124 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_137 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_123 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _rmask_T_138 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_140 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_142 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_144 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_146 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_148 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_150 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_152 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_154 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_156 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_158 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_160 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_162 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] rmask_3 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rData_T_19 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5890 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire [31:0] _GEN_5891 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5892 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [31:0] rData_3 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5893 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _T_1095 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _T_1096 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _T_1097 = ~_T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:63]
  wire [31:0] _T_1098 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mepc_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mepc_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire  _T_1075 = csrAddr == 12'h341; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _next_csr_mepc_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mepc_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire  _T_1051 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_1052 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _T_1053 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _rData_T_14 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _rData_T_15 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _rData_T_16 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _rData_T_17 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire  _has_T_323 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_321 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_319 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_317 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_315 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_313 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_311 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_309 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_307 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_305 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_303 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_301 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_299 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_297 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_298 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_300 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_302 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_304 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_306 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_308 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_310 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_312 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_314 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_316 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_318 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_320 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_322 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  has_11 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _nowCSR_T_80 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_78 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_76 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_74 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_72 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_70 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_68 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_66 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_64 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_62 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_60 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_58 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_56 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_54 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_55 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_57 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_59 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_61 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_63 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_65 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_67 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_69 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_71 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_73 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_75 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_77 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_79 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] nowCSR_2 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _rData_T_12 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _rmask_T_122 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_95 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_120 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_94 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_118 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_93 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_116 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_92 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_114 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_91 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_112 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_90 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_110 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_89 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_108 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_88 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_106 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_87 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_104 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_86 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_102 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_85 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_100 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_84 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_98 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_83 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_96 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_82 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _rmask_T_97 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_99 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_101 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_103 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_105 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_107 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_109 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_111 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_113 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_115 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_117 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_119 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_121 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] rmask_2 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rData_T_13 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5718 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire [31:0] _GEN_5719 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5720 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [31:0] rData_2 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5721 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _T_1055 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _T_1056 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _T_1057 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mepc_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mepc_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire  _T_1034 = csrAddr == 12'h341; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _next_csr_mepc_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mepc_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _T_1016 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mepc_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mepc_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  _T_1000 = csrAddr == 12'h341; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _next_csr_mepc_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mepc_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire  _T_976 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_977 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _T_978 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _rData_T_8 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _rData_T_9 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _rData_T_10 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _rData_T_11 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire  _has_T_188 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_186 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_184 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_182 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_180 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_178 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_176 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_174 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_172 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_170 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_168 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_166 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_164 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_162 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_163 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_165 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_167 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_169 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_171 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_173 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_175 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_177 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_179 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_181 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_183 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_185 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_187 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  has_6 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _nowCSR_T_53 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_51 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_49 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_47 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_45 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_43 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_41 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_39 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_37 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_35 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_33 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_31 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_29 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_27 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_28 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_30 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_32 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_34 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_36 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_38 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_40 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_42 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_44 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_46 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_48 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_50 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_52 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] nowCSR_1 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _rData_T_6 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _rmask_T_81 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_54 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_79 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_53 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_77 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_52 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_75 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_51 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_73 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_50 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_71 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_49 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_69 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_48 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_67 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_47 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_65 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_46 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_63 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_45 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_61 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_44 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_59 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_43 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_57 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_42 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_55 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_41 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _rmask_T_56 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_58 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_60 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_62 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_64 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_66 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_68 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_70 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_72 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_74 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_76 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_78 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_80 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] rmask_1 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rData_T_7 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5358 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire [31:0] _GEN_5359 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5360 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [31:0] rData_1 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5361 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _T_980 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _now_reg_rs1_73 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _T_981 = ~_GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:63]
  wire [31:0] _T_982 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mepc_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mepc_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire  _T_960 = csrAddr == 12'h341; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _next_csr_mepc_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mepc_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire  _T_937 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_938 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _T_939 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _rData_T_2 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _rData_T_3 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _rData_T_4 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _rData_T_5 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire  _has_T_107 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_105 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_103 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_101 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_99 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_97 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_95 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_93 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_91 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_89 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_87 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_85 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_83 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_81 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_82 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_84 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_86 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_88 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_90 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_92 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_94 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_96 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_98 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_100 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_102 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_104 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _has_T_106 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  has_3 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _nowCSR_T_26 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_24 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_22 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_20 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_18 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_16 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_14 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_12 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_10 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_8 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_6 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_4 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T_2 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _nowCSR_T = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_1 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_3 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_5 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_7 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_9 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_11 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_13 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_15 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_17 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_19 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_21 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_23 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _nowCSR_T_25 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] nowCSR = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _rData_T = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _rmask_T_40 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_13 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_38 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_36 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_11 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_34 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_10 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_32 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_30 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_8 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_28 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_7 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_26 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_24 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_5 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_22 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_4 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_20 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_18 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_2 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_16 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_1 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _rmask_T_14 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _rmask_T_15 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_17 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_19 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_21 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_23 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_25 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_27 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_29 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_31 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_33 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_35 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_37 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rmask_T_39 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] rmask = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _rData_T_1 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5186 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire [31:0] _GEN_5187 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5188 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [31:0] rData = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5189 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _T_941 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _now_reg_rs1_72 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _T_942 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mepc_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mepc_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire  _T_920 = csrAddr == 12'h341; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _next_csr_mepc_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mepc_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _now_reg_rs1_68 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mepc_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mepc_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mepc_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5037 = csrAddr == 12'h341 ? _GEN_31 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5047 = has_15 ? _GEN_5037 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5091 = _T_1089 ? _GEN_5047 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5145 = _T_894 ? _GEN_5091 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5197 = csrAddr == 12'h341 ? _T_942 : _GEN_5145; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5207 = has_15 ? _GEN_5197 : _GEN_5145; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5219 = _T_1090 ? _GEN_5207 : _GEN_5145; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5263 = _T_1049 ? _GEN_5219 : _GEN_5145; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5317 = _T_927 ? _GEN_5263 : _GEN_5145; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5369 = csrAddr == 12'h341 ? _T_982 : _GEN_5317; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5379 = has_15 ? _GEN_5369 : _GEN_5317; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5391 = _T_1090 ? _GEN_5379 : _GEN_5317; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5435 = _T_1089 ? _GEN_5391 : _GEN_5317; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5489 = _T_967 ? _GEN_5435 : _GEN_5317; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5569 = csrAddr == 12'h341 ? _T_1096 : _GEN_5489; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5579 = has_15 ? _GEN_5569 : _GEN_5489; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5623 = _T_1089 ? _GEN_5579 : _GEN_5489; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5677 = _T_1007 ? _GEN_5623 : _GEN_5489; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5729 = csrAddr == 12'h341 ? _T_1057 : _GEN_5677; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5739 = has_15 ? _GEN_5729 : _GEN_5677; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5751 = _T_1090 ? _GEN_5739 : _GEN_5677; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5795 = ~isIllegalWrite_4 ? _GEN_5751 : _GEN_5677; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5849 = _T_1041 ? _GEN_5795 : _GEN_5677; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5901 = csrAddr == 12'h341 ? _T_1098 : _GEN_5849; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5911 = has_15 ? _GEN_5901 : _GEN_5849; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5923 = rs1 != 5'h0 ? _GEN_5911 : _GEN_5849; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5967 = ~isIllegalWrite_5 ? _GEN_5923 : _GEN_5849; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_6021 = _T_1082 ? _GEN_5967 : _GEN_5849; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire  _T_1141 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_6061 = _T_1123 ? io_now_pc : _GEN_6021; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 186:35]
  wire [31:0] _GEN_6085 = delegS ? _GEN_6021 : _GEN_6061; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [31:0] _GEN_6099 = raiseExceptionIntr ? _GEN_6085 : _GEN_6021; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_mepc = io_valid ? _GEN_6099 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6198 = next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _retTarget_T_1 = next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [1:0] _mstatusOld_WIRE_2_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_31 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _GEN_4925 = io_now_internal_privilegeMode == 2'h3 ? mstatusOld_mpp : _GEN_4920; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 92:35]
  wire [31:0] _GEN_4926 = io_now_internal_privilegeMode == 2'h3 ? _next_csr_mstatus_T_1 : _GEN_4921; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:24 88:48]
  wire [31:0] _GEN_4927 = io_now_internal_privilegeMode == 2'h3 ? next_csr_mepc : next_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 101:24 88:48]
  wire  _GEN_4928 = io_now_internal_privilegeMode == 2'h3 | _GEN_4923; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 103:25 88:48]
  wire [31:0] _GEN_4929 = io_now_internal_privilegeMode == 2'h3 ? io_now_csr_mepc : _GEN_4924; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 104:25 88:48]
  wire [2:0] _GEN_4935 = _T_875 ? inst[14:12] : _GEN_4914; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4937 = _T_875 ? inst[6:0] : _GEN_4916; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [1:0] _GEN_4939 = _T_875 ? _GEN_4925 : _GEN_4920; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _GEN_4940 = _T_875 ? _GEN_4926 : _GEN_4921; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] retTarget = _T_875 ? _GEN_4927 : next_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_4942 = _T_875 ? _GEN_4928 : _GEN_4923; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _GEN_4943 = _T_875 ? _GEN_4929 : _GEN_4924; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [2:0] _funct3_T_65 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_886 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_4949 = _T_882 ? inst[14:12] : _GEN_4935; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4951 = _T_882 ? inst[6:0] : _GEN_4937; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [2:0] _funct3_T_66 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_892 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_4956 = _T_888 ? inst[14:12] : _GEN_4949; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_4958 = _T_888 ? inst[6:0] : _GEN_4951; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [2:0] _funct3_T_67 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_898 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _T_902 = rd != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:17]
  wire  _next_reg_has_T = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_1 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_2 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_3 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_4 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_5 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_6 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_7 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_8 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_9 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_10 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_11 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_12 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_13 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_14 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_15 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_16 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_17 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_18 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_19 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_20 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_21 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_22 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_23 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_24 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_25 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_26 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  next_reg_has = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_nowCSR_T = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_1 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_2 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_3 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_4 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_5 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_6 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_7 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_8 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_9 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_10 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_11 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_12 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_13 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_14 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_15 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_16 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_17 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_18 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_19 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_20 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_21 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_22 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_23 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_24 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_25 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_26 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] next_reg_nowCSR = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rmask_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_1 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_2 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_4 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_5 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_7 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_8 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_10 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_11 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_13 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _next_reg_rmask_T_14 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_15 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_16 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_17 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_18 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_19 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_20 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_21 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_22 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_23 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_24 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_25 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_26 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_27 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_28 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_29 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_30 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_31 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_32 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_33 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_34 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_35 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_36 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_37 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_38 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_39 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_40 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] next_reg_rmask = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_T_181 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] _next_reg_rData_T = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rData_T_1 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_4962 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire  _next_reg_T_182 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_183 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _next_reg_rData_T_2 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _next_reg_rData_T_3 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _next_reg_rData_T_4 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _next_reg_rData_T_5 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [31:0] _GEN_4963 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_4964 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_184 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] next_reg_rData = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_4965 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_T_185 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_rd_42 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_4966 = 5'h0 == rd ? rData_3 : _GEN_4868; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4967 = 5'h1 == rd ? rData_3 : _GEN_4869; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4968 = 5'h2 == rd ? rData_3 : _GEN_4870; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4969 = 5'h3 == rd ? rData_3 : _GEN_4871; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4970 = 5'h4 == rd ? rData_3 : _GEN_4872; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4971 = 5'h5 == rd ? rData_3 : _GEN_4873; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4972 = 5'h6 == rd ? rData_3 : _GEN_4874; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4973 = 5'h7 == rd ? rData_3 : _GEN_4875; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4974 = 5'h8 == rd ? rData_3 : _GEN_4876; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4975 = 5'h9 == rd ? rData_3 : _GEN_4877; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4976 = 5'ha == rd ? rData_3 : _GEN_4878; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4977 = 5'hb == rd ? rData_3 : _GEN_4879; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4978 = 5'hc == rd ? rData_3 : _GEN_4880; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4979 = 5'hd == rd ? rData_3 : _GEN_4881; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4980 = 5'he == rd ? rData_3 : _GEN_4882; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4981 = 5'hf == rd ? rData_3 : _GEN_4883; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4982 = 5'h10 == rd ? rData_3 : _GEN_4884; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4983 = 5'h11 == rd ? rData_3 : _GEN_4885; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4984 = 5'h12 == rd ? rData_3 : _GEN_4886; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4985 = 5'h13 == rd ? rData_3 : _GEN_4887; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4986 = 5'h14 == rd ? rData_3 : _GEN_4888; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4987 = 5'h15 == rd ? rData_3 : _GEN_4889; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4988 = 5'h16 == rd ? rData_3 : _GEN_4890; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4989 = 5'h17 == rd ? rData_3 : _GEN_4891; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4990 = 5'h18 == rd ? rData_3 : _GEN_4892; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4991 = 5'h19 == rd ? rData_3 : _GEN_4893; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4992 = 5'h1a == rd ? rData_3 : _GEN_4894; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4993 = 5'h1b == rd ? rData_3 : _GEN_4895; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4994 = 5'h1c == rd ? rData_3 : _GEN_4896; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4995 = 5'h1d == rd ? rData_3 : _GEN_4897; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4996 = 5'h1e == rd ? rData_3 : _GEN_4898; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4997 = 5'h1f == rd ? rData_3 : _GEN_4899; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [31:0] _GEN_4998 = rd != 5'h0 ? _GEN_4966 : _GEN_4868; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_4999 = rd != 5'h0 ? _GEN_4967 : _GEN_4869; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5000 = rd != 5'h0 ? _GEN_4968 : _GEN_4870; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5001 = rd != 5'h0 ? _GEN_4969 : _GEN_4871; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5002 = rd != 5'h0 ? _GEN_4970 : _GEN_4872; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5003 = rd != 5'h0 ? _GEN_4971 : _GEN_4873; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5004 = rd != 5'h0 ? _GEN_4972 : _GEN_4874; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5005 = rd != 5'h0 ? _GEN_4973 : _GEN_4875; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5006 = rd != 5'h0 ? _GEN_4974 : _GEN_4876; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5007 = rd != 5'h0 ? _GEN_4975 : _GEN_4877; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5008 = rd != 5'h0 ? _GEN_4976 : _GEN_4878; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5009 = rd != 5'h0 ? _GEN_4977 : _GEN_4879; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5010 = rd != 5'h0 ? _GEN_4978 : _GEN_4880; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5011 = rd != 5'h0 ? _GEN_4979 : _GEN_4881; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5012 = rd != 5'h0 ? _GEN_4980 : _GEN_4882; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5013 = rd != 5'h0 ? _GEN_4981 : _GEN_4883; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5014 = rd != 5'h0 ? _GEN_4982 : _GEN_4884; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5015 = rd != 5'h0 ? _GEN_4983 : _GEN_4885; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5016 = rd != 5'h0 ? _GEN_4984 : _GEN_4886; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5017 = rd != 5'h0 ? _GEN_4985 : _GEN_4887; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5018 = rd != 5'h0 ? _GEN_4986 : _GEN_4888; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5019 = rd != 5'h0 ? _GEN_4987 : _GEN_4889; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5020 = rd != 5'h0 ? _GEN_4988 : _GEN_4890; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5021 = rd != 5'h0 ? _GEN_4989 : _GEN_4891; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5022 = rd != 5'h0 ? _GEN_4990 : _GEN_4892; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5023 = rd != 5'h0 ? _GEN_4991 : _GEN_4893; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5024 = rd != 5'h0 ? _GEN_4992 : _GEN_4894; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5025 = rd != 5'h0 ? _GEN_4993 : _GEN_4895; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5026 = rd != 5'h0 ? _GEN_4994 : _GEN_4896; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5027 = rd != 5'h0 ? _GEN_4995 : _GEN_4897; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5028 = rd != 5'h0 ? _GEN_4996 : _GEN_4898; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [31:0] _GEN_5029 = rd != 5'h0 ? _GEN_4997 : _GEN_4899; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire  _T_903 = csrAddr == 12'h301; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_904 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_misa_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_misa_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_61 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_misa_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_misa_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5030 = csrAddr == 12'h301 ? _GEN_31 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_905 = csrAddr == 12'hf11; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_906 = csrAddr == 12'hf12; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_907 = csrAddr == 12'hf13; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_908 = csrAddr == 12'hf14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_909 = csrAddr == 12'h300; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_910 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_2 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mstatus_T_4 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mstatus_T_5 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_62 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mstatus_T_6 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mstatus_T_7 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mstatus_mstatusOld_WIRE_1 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  next_csr_mstatus_mstatusOld_pad4 = _GEN_31[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sie = _GEN_31[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_pad3 = _GEN_31[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mie = _GEN_31[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_pad2 = _GEN_31[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_spie = _GEN_31[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_ube = _GEN_31[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mpie = _GEN_31[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_spp = _GEN_31[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_vs = _GEN_31[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_mpp = _GEN_31[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_fs = _GEN_31[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_xs = _GEN_31[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mprv = _GEN_31[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sum = _GEN_31[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mxr = _GEN_31[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_tvm = _GEN_31[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_tw = _GEN_31[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_tsr = _GEN_31[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] next_csr_mstatus_mstatusOld_pad0 = _GEN_31[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sd = _GEN_31[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_fs = next_csr_mstatus_mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_11 = next_csr_mstatus_mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusNew_T = next_csr_mstatus_mstatusOld_fs == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:42]
  wire  _next_csr_mstatus_mstatusOld_WIRE_sie = next_csr_mstatus_mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_1 = next_csr_mstatus_mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_pad4 = next_csr_mstatus_mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T = next_csr_mstatus_mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_lo = {next_csr_mstatus_mstatusOld_sie,next_csr_mstatus_mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_pad2 = next_csr_mstatus_mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_4 = next_csr_mstatus_mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_mie = next_csr_mstatus_mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_3 = next_csr_mstatus_mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_hi_hi = {next_csr_mstatus_mstatusOld_pad2,next_csr_mstatus_mstatusOld_mie
    }; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_pad3 = next_csr_mstatus_mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_2 = next_csr_mstatus_mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_lo_hi = {next_csr_mstatus_mstatusOld_pad2,next_csr_mstatus_mstatusOld_mie,
    next_csr_mstatus_mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [4:0] next_csr_mstatus_mstatusNew_lo_lo = {next_csr_mstatus_mstatusOld_pad2,next_csr_mstatus_mstatusOld_mie,
    next_csr_mstatus_mstatusOld_pad3,next_csr_mstatus_mstatusOld_sie,next_csr_mstatus_mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_ube = next_csr_mstatus_mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_6 = next_csr_mstatus_mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_spie = next_csr_mstatus_mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_5 = next_csr_mstatus_mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_hi_lo = {next_csr_mstatus_mstatusOld_ube,next_csr_mstatus_mstatusOld_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_vs = next_csr_mstatus_mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_9 = next_csr_mstatus_mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_spp = next_csr_mstatus_mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_8 = next_csr_mstatus_mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_hi_hi_hi = {next_csr_mstatus_mstatusOld_vs,next_csr_mstatus_mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_mpie = next_csr_mstatus_mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_7 = next_csr_mstatus_mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_lo_hi_hi = {next_csr_mstatus_mstatusOld_vs,next_csr_mstatus_mstatusOld_spp,
    next_csr_mstatus_mstatusOld_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_hi = {next_csr_mstatus_mstatusOld_vs,next_csr_mstatus_mstatusOld_spp,
    next_csr_mstatus_mstatusOld_mpie,next_csr_mstatus_mstatusOld_ube,next_csr_mstatus_mstatusOld_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [10:0] next_csr_mstatus_mstatusNew_lo = {next_csr_mstatus_mstatusOld_vs,next_csr_mstatus_mstatusOld_spp,
    next_csr_mstatus_mstatusOld_mpie,next_csr_mstatus_mstatusOld_ube,next_csr_mstatus_mstatusOld_spie,
    next_csr_mstatus_mstatusOld_pad2,next_csr_mstatus_mstatusOld_mie,next_csr_mstatus_mstatusOld_pad3,
    next_csr_mstatus_mstatusOld_sie,next_csr_mstatus_mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_mpp = next_csr_mstatus_mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_10 = next_csr_mstatus_mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_lo = {next_csr_mstatus_mstatusOld_fs,next_csr_mstatus_mstatusOld_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_sum = next_csr_mstatus_mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_14 = next_csr_mstatus_mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_mprv = next_csr_mstatus_mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_13 = next_csr_mstatus_mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_lo_hi_hi = {next_csr_mstatus_mstatusOld_sum,next_csr_mstatus_mstatusOld_mprv
    }; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_xs = next_csr_mstatus_mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_12 = next_csr_mstatus_mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_hi = {next_csr_mstatus_mstatusOld_sum,next_csr_mstatus_mstatusOld_mprv,
    next_csr_mstatus_mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [7:0] next_csr_mstatus_mstatusNew_hi_lo = {next_csr_mstatus_mstatusOld_sum,next_csr_mstatus_mstatusOld_mprv,
    next_csr_mstatus_mstatusOld_xs,next_csr_mstatus_mstatusOld_fs,next_csr_mstatus_mstatusOld_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_tw = next_csr_mstatus_mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_17 = next_csr_mstatus_mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_tvm = next_csr_mstatus_mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_16 = next_csr_mstatus_mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_hi_lo_hi = {next_csr_mstatus_mstatusOld_tw,next_csr_mstatus_mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_mxr = next_csr_mstatus_mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_15 = next_csr_mstatus_mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_hi_hi_lo = {next_csr_mstatus_mstatusOld_tw,next_csr_mstatus_mstatusOld_tvm,
    next_csr_mstatus_mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_sd = next_csr_mstatus_mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_20 = next_csr_mstatus_mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_WIRE_pad0 = next_csr_mstatus_mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_T_19 = next_csr_mstatus_mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusNew_hi_hi_hi_hi = {next_csr_mstatus_mstatusOld_sd,next_csr_mstatus_mstatusOld_pad0}
    ; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_tsr = next_csr_mstatus_mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_18 = next_csr_mstatus_mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [9:0] next_csr_mstatus_mstatusNew_hi_hi_hi = {next_csr_mstatus_mstatusOld_sd,next_csr_mstatus_mstatusOld_pad0,
    next_csr_mstatus_mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [12:0] next_csr_mstatus_mstatusNew_hi_hi = {next_csr_mstatus_mstatusOld_sd,next_csr_mstatus_mstatusOld_pad0,
    next_csr_mstatus_mstatusOld_tsr,next_csr_mstatus_mstatusOld_tw,next_csr_mstatus_mstatusOld_tvm,
    next_csr_mstatus_mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [20:0] next_csr_mstatus_mstatusNew_hi = {next_csr_mstatus_mstatusOld_sd,next_csr_mstatus_mstatusOld_pad0,
    next_csr_mstatus_mstatusOld_tsr,next_csr_mstatus_mstatusOld_tw,next_csr_mstatus_mstatusOld_tvm,
    next_csr_mstatus_mstatusOld_mxr,next_csr_mstatus_mstatusNew_hi_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [31:0] _next_csr_mstatus_mstatusNew_T_1 = {next_csr_mstatus_mstatusOld_sd,next_csr_mstatus_mstatusOld_pad0,
    next_csr_mstatus_mstatusOld_tsr,next_csr_mstatus_mstatusOld_tw,next_csr_mstatus_mstatusOld_tvm,
    next_csr_mstatus_mstatusOld_mxr,next_csr_mstatus_mstatusNew_hi_lo,next_csr_mstatus_mstatusNew_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [30:0] _next_csr_mstatus_mstatusNew_T_2 = _next_csr_mstatus_mstatusNew_T_1[30:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:72]
  wire [31:0] next_csr_mstatus_mstatusNew = {next_csr_mstatus_mstatusOld_fs == 2'h3,_next_csr_mstatus_mstatusNew_T_1[30:
    0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [31:0] _GEN_5031 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew : _GEN_4940; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_911 = csrAddr == 12'h340; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_912 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mscratch_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mscratch_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_63 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mscratch_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mscratch_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5032 = csrAddr == 12'h340 ? _GEN_31 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_913 = csrAddr == 12'h305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_914 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtvec_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtvec_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_64 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mtvec_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mtvec_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5033 = csrAddr == 12'h305 ? _GEN_31 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_915 = csrAddr == 12'h306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_916 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcounteren_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcounteren_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_65 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mcounteren_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mcounteren_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5034 = csrAddr == 12'h306 ? _GEN_31 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_917 = csrAddr == 12'h344; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [10:0] _next_csr_mip_T = 11'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mip_T_1 = io_now_csr_mip & 32'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _now_reg_rs1_66 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mip_T_2 = _GEN_31 & 32'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [31:0] _next_csr_mip_T_3 = _next_csr_mip_T_1 | _next_csr_mip_T_2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [31:0] _GEN_5035 = csrAddr == 12'h344 ? _next_csr_mip_T_3 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_918 = csrAddr == 12'h304; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_919 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mie_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mie_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_67 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mie_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mie_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5036 = csrAddr == 12'h304 ? _GEN_31 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _T_921 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire  _T_922 = csrAddr == 12'h342; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_923 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcause_T_2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcause_T_3 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_69 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mcause_T_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mcause_T_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5038 = csrAddr == 12'h342 ? _GEN_31 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_924 = csrAddr == 12'h343; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_925 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtval_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtval_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _now_reg_rs1_70 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mtval_T_22 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_csr_mtval_T_23 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5039 = csrAddr == 12'h343 ? _GEN_31 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5040 = has_15 ? _GEN_5030 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5041 = has_15 ? _GEN_5031 : _GEN_4940; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5042 = has_15 ? _GEN_5032 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5043 = has_15 ? _GEN_5033 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5044 = has_15 ? _GEN_5034 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5045 = has_15 ? _GEN_5035 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5046 = has_15 ? _GEN_5036 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5048 = has_15 ? _GEN_5038 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_5049 = has_15 ? _GEN_5039 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5052 = _T_1089 ? _GEN_4998 : _GEN_4868; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5053 = _T_1089 ? _GEN_4999 : _GEN_4869; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5054 = _T_1089 ? _GEN_5000 : _GEN_4870; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5055 = _T_1089 ? _GEN_5001 : _GEN_4871; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5056 = _T_1089 ? _GEN_5002 : _GEN_4872; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5057 = _T_1089 ? _GEN_5003 : _GEN_4873; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5058 = _T_1089 ? _GEN_5004 : _GEN_4874; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5059 = _T_1089 ? _GEN_5005 : _GEN_4875; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5060 = _T_1089 ? _GEN_5006 : _GEN_4876; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5061 = _T_1089 ? _GEN_5007 : _GEN_4877; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5062 = _T_1089 ? _GEN_5008 : _GEN_4878; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5063 = _T_1089 ? _GEN_5009 : _GEN_4879; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5064 = _T_1089 ? _GEN_5010 : _GEN_4880; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5065 = _T_1089 ? _GEN_5011 : _GEN_4881; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5066 = _T_1089 ? _GEN_5012 : _GEN_4882; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5067 = _T_1089 ? _GEN_5013 : _GEN_4883; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5068 = _T_1089 ? _GEN_5014 : _GEN_4884; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5069 = _T_1089 ? _GEN_5015 : _GEN_4885; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5070 = _T_1089 ? _GEN_5016 : _GEN_4886; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5071 = _T_1089 ? _GEN_5017 : _GEN_4887; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5072 = _T_1089 ? _GEN_5018 : _GEN_4888; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5073 = _T_1089 ? _GEN_5019 : _GEN_4889; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5074 = _T_1089 ? _GEN_5020 : _GEN_4890; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5075 = _T_1089 ? _GEN_5021 : _GEN_4891; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5076 = _T_1089 ? _GEN_5022 : _GEN_4892; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5077 = _T_1089 ? _GEN_5023 : _GEN_4893; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5078 = _T_1089 ? _GEN_5024 : _GEN_4894; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5079 = _T_1089 ? _GEN_5025 : _GEN_4895; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5080 = _T_1089 ? _GEN_5026 : _GEN_4896; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5081 = _T_1089 ? _GEN_5027 : _GEN_4897; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5082 = _T_1089 ? _GEN_5028 : _GEN_4898; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5083 = _T_1089 ? _GEN_5029 : _GEN_4899; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5084 = _T_1089 ? _GEN_5040 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5085 = _T_1089 ? _GEN_5041 : _GEN_4940; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5086 = _T_1089 ? _GEN_5042 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5087 = _T_1089 ? _GEN_5043 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5088 = _T_1089 ? _GEN_5044 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5089 = _T_1089 ? _GEN_5045 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5090 = _T_1089 ? _GEN_5046 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5092 = _T_1089 ? _GEN_5048 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [31:0] _GEN_5093 = _T_1089 ? _GEN_5049 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [2:0] _GEN_5099 = _T_894 ? inst[14:12] : _GEN_4956; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5101 = _T_894 ? inst[6:0] : _GEN_4958; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_5106 = _T_894 ? _GEN_5052 : _GEN_4868; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5107 = _T_894 ? _GEN_5053 : _GEN_4869; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5108 = _T_894 ? _GEN_5054 : _GEN_4870; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5109 = _T_894 ? _GEN_5055 : _GEN_4871; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5110 = _T_894 ? _GEN_5056 : _GEN_4872; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5111 = _T_894 ? _GEN_5057 : _GEN_4873; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5112 = _T_894 ? _GEN_5058 : _GEN_4874; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5113 = _T_894 ? _GEN_5059 : _GEN_4875; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5114 = _T_894 ? _GEN_5060 : _GEN_4876; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5115 = _T_894 ? _GEN_5061 : _GEN_4877; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5116 = _T_894 ? _GEN_5062 : _GEN_4878; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5117 = _T_894 ? _GEN_5063 : _GEN_4879; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5118 = _T_894 ? _GEN_5064 : _GEN_4880; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5119 = _T_894 ? _GEN_5065 : _GEN_4881; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5120 = _T_894 ? _GEN_5066 : _GEN_4882; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5121 = _T_894 ? _GEN_5067 : _GEN_4883; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5122 = _T_894 ? _GEN_5068 : _GEN_4884; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5123 = _T_894 ? _GEN_5069 : _GEN_4885; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5124 = _T_894 ? _GEN_5070 : _GEN_4886; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5125 = _T_894 ? _GEN_5071 : _GEN_4887; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5126 = _T_894 ? _GEN_5072 : _GEN_4888; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5127 = _T_894 ? _GEN_5073 : _GEN_4889; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5128 = _T_894 ? _GEN_5074 : _GEN_4890; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5129 = _T_894 ? _GEN_5075 : _GEN_4891; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5130 = _T_894 ? _GEN_5076 : _GEN_4892; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5131 = _T_894 ? _GEN_5077 : _GEN_4893; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5132 = _T_894 ? _GEN_5078 : _GEN_4894; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5133 = _T_894 ? _GEN_5079 : _GEN_4895; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5134 = _T_894 ? _GEN_5080 : _GEN_4896; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5135 = _T_894 ? _GEN_5081 : _GEN_4897; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5136 = _T_894 ? _GEN_5082 : _GEN_4898; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5137 = _T_894 ? _GEN_5083 : _GEN_4899; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5138 = _T_894 ? _GEN_5084 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5139 = _T_894 ? _GEN_5085 : _GEN_4940; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5140 = _T_894 ? _GEN_5086 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5141 = _T_894 ? _GEN_5087 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5142 = _T_894 ? _GEN_5088 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5143 = _T_894 ? _GEN_5089 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5144 = _T_894 ? _GEN_5090 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5146 = _T_894 ? _GEN_5092 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [31:0] _GEN_5147 = _T_894 ? _GEN_5093 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [2:0] _funct3_T_68 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_931 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _next_reg_has_T_27 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_28 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_29 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_30 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_31 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_32 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_33 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_34 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_35 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_36 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_37 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_38 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_39 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_40 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_41 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_42 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_43 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_44 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_45 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_46 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_47 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_48 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_49 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_50 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_51 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_52 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_53 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  next_reg_has_1 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_nowCSR_T_27 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_28 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_29 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_30 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_31 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_32 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_33 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_34 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_35 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_36 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_37 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_38 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_39 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_40 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_41 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_42 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_43 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_44 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_45 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_46 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_47 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_48 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_49 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_50 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_51 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_52 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_53 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] next_reg_nowCSR_1 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rmask_T_41 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_42 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_43 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_44 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_45 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_46 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_47 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_48 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_49 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_50 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_51 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_52 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_53 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_54 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _next_reg_rmask_T_55 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_56 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_57 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_58 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_59 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_60 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_61 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_62 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_63 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_64 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_65 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_66 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_67 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_68 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_69 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_70 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_71 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_72 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_73 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_74 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_75 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_76 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_77 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_78 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_79 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_80 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_81 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] next_reg_rmask_1 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_T_186 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] _next_reg_rData_T_6 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rData_T_7 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5150 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire  _next_reg_T_187 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_188 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _next_reg_rData_T_8 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _next_reg_rData_T_9 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _next_reg_rData_T_10 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _next_reg_rData_T_11 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [31:0] _GEN_5151 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5152 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_189 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] next_reg_rData_1 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5153 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_T_190 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_rd_43 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5154 = 5'h0 == rd ? rData_3 : _GEN_5106; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5155 = 5'h1 == rd ? rData_3 : _GEN_5107; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5156 = 5'h2 == rd ? rData_3 : _GEN_5108; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5157 = 5'h3 == rd ? rData_3 : _GEN_5109; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5158 = 5'h4 == rd ? rData_3 : _GEN_5110; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5159 = 5'h5 == rd ? rData_3 : _GEN_5111; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5160 = 5'h6 == rd ? rData_3 : _GEN_5112; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5161 = 5'h7 == rd ? rData_3 : _GEN_5113; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5162 = 5'h8 == rd ? rData_3 : _GEN_5114; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5163 = 5'h9 == rd ? rData_3 : _GEN_5115; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5164 = 5'ha == rd ? rData_3 : _GEN_5116; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5165 = 5'hb == rd ? rData_3 : _GEN_5117; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5166 = 5'hc == rd ? rData_3 : _GEN_5118; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5167 = 5'hd == rd ? rData_3 : _GEN_5119; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5168 = 5'he == rd ? rData_3 : _GEN_5120; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5169 = 5'hf == rd ? rData_3 : _GEN_5121; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5170 = 5'h10 == rd ? rData_3 : _GEN_5122; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5171 = 5'h11 == rd ? rData_3 : _GEN_5123; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5172 = 5'h12 == rd ? rData_3 : _GEN_5124; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5173 = 5'h13 == rd ? rData_3 : _GEN_5125; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5174 = 5'h14 == rd ? rData_3 : _GEN_5126; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5175 = 5'h15 == rd ? rData_3 : _GEN_5127; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5176 = 5'h16 == rd ? rData_3 : _GEN_5128; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5177 = 5'h17 == rd ? rData_3 : _GEN_5129; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5178 = 5'h18 == rd ? rData_3 : _GEN_5130; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5179 = 5'h19 == rd ? rData_3 : _GEN_5131; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5180 = 5'h1a == rd ? rData_3 : _GEN_5132; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5181 = 5'h1b == rd ? rData_3 : _GEN_5133; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5182 = 5'h1c == rd ? rData_3 : _GEN_5134; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5183 = 5'h1d == rd ? rData_3 : _GEN_5135; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5184 = 5'h1e == rd ? rData_3 : _GEN_5136; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [31:0] _GEN_5185 = 5'h1f == rd ? rData_3 : _GEN_5137; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire  _T_940 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_943 = csrAddr == 12'h301; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_944 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_misa_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_misa_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_misa_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5190 = csrAddr == 12'h301 ? _T_942 : _GEN_5138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_945 = csrAddr == 12'hf11; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_946 = csrAddr == 12'hf12; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_947 = csrAddr == 12'hf13; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_948 = csrAddr == 12'hf14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_949 = csrAddr == 12'h300; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_950 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_8 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_9 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mstatus_T_10 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mstatus_T_11 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_12 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mstatus_T_13 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mstatus_mstatusOld_WIRE_3 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire  next_csr_mstatus_mstatusOld_1_pad4 = _T_942[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sie = _T_942[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_pad3 = _T_942[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mie = _T_942[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_pad2 = _T_942[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_spie = _T_942[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_ube = _T_942[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mpie = _T_942[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_spp = _T_942[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_vs = _T_942[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_mpp = _T_942[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_fs = _T_942[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_xs = _T_942[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mprv = _T_942[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sum = _T_942[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mxr = _T_942[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_tvm = _T_942[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_tw = _T_942[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_tsr = _T_942[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] next_csr_mstatus_mstatusOld_1_pad0 = _T_942[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sd = _T_942[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_2_fs = next_csr_mstatus_mstatusOld_1_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_32 = next_csr_mstatus_mstatusOld_1_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusNew_T_3 = next_csr_mstatus_mstatusOld_1_fs == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:42]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_sie = next_csr_mstatus_mstatusOld_1_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_22 = next_csr_mstatus_mstatusOld_1_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_pad4 = next_csr_mstatus_mstatusOld_1_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_21 = next_csr_mstatus_mstatusOld_1_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_lo_1 = {next_csr_mstatus_mstatusOld_1_sie,
    next_csr_mstatus_mstatusOld_1_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_pad2 = next_csr_mstatus_mstatusOld_1_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_25 = next_csr_mstatus_mstatusOld_1_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_mie = next_csr_mstatus_mstatusOld_1_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_24 = next_csr_mstatus_mstatusOld_1_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_pad2,
    next_csr_mstatus_mstatusOld_1_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_pad3 = next_csr_mstatus_mstatusOld_1_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_23 = next_csr_mstatus_mstatusOld_1_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_lo_hi_1 = {next_csr_mstatus_mstatusOld_1_pad2,
    next_csr_mstatus_mstatusOld_1_mie,next_csr_mstatus_mstatusOld_1_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [4:0] next_csr_mstatus_mstatusNew_lo_lo_1 = {next_csr_mstatus_mstatusOld_1_pad2,next_csr_mstatus_mstatusOld_1_mie
    ,next_csr_mstatus_mstatusOld_1_pad3,next_csr_mstatus_mstatusOld_1_sie,next_csr_mstatus_mstatusOld_1_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_ube = next_csr_mstatus_mstatusOld_1_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_27 = next_csr_mstatus_mstatusOld_1_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_spie = next_csr_mstatus_mstatusOld_1_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_26 = next_csr_mstatus_mstatusOld_1_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_hi_lo_1 = {next_csr_mstatus_mstatusOld_1_ube,
    next_csr_mstatus_mstatusOld_1_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_2_vs = next_csr_mstatus_mstatusOld_1_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_30 = next_csr_mstatus_mstatusOld_1_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_spp = next_csr_mstatus_mstatusOld_1_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_29 = next_csr_mstatus_mstatusOld_1_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_hi_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_vs,
    next_csr_mstatus_mstatusOld_1_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_mpie = next_csr_mstatus_mstatusOld_1_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_28 = next_csr_mstatus_mstatusOld_1_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_lo_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_vs,
    next_csr_mstatus_mstatusOld_1_spp,next_csr_mstatus_mstatusOld_1_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_hi_1 = {next_csr_mstatus_mstatusOld_1_vs,next_csr_mstatus_mstatusOld_1_spp,
    next_csr_mstatus_mstatusOld_1_mpie,next_csr_mstatus_mstatusOld_1_ube,next_csr_mstatus_mstatusOld_1_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [10:0] next_csr_mstatus_mstatusNew_lo_1 = {next_csr_mstatus_mstatusOld_1_vs,next_csr_mstatus_mstatusOld_1_spp,
    next_csr_mstatus_mstatusOld_1_mpie,next_csr_mstatus_mstatusOld_1_ube,next_csr_mstatus_mstatusOld_1_spie,
    next_csr_mstatus_mstatusOld_1_pad2,next_csr_mstatus_mstatusOld_1_mie,next_csr_mstatus_mstatusOld_1_pad3,
    next_csr_mstatus_mstatusOld_1_sie,next_csr_mstatus_mstatusOld_1_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_2_mpp = next_csr_mstatus_mstatusOld_1_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_31 = next_csr_mstatus_mstatusOld_1_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_lo_1 = {next_csr_mstatus_mstatusOld_1_fs,
    next_csr_mstatus_mstatusOld_1_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_sum = next_csr_mstatus_mstatusOld_1_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_35 = next_csr_mstatus_mstatusOld_1_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_mprv = next_csr_mstatus_mstatusOld_1_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_34 = next_csr_mstatus_mstatusOld_1_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_lo_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_sum,
    next_csr_mstatus_mstatusOld_1_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_2_xs = next_csr_mstatus_mstatusOld_1_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_33 = next_csr_mstatus_mstatusOld_1_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_hi_1 = {next_csr_mstatus_mstatusOld_1_sum,
    next_csr_mstatus_mstatusOld_1_mprv,next_csr_mstatus_mstatusOld_1_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [7:0] next_csr_mstatus_mstatusNew_hi_lo_1 = {next_csr_mstatus_mstatusOld_1_sum,next_csr_mstatus_mstatusOld_1_mprv
    ,next_csr_mstatus_mstatusOld_1_xs,next_csr_mstatus_mstatusOld_1_fs,next_csr_mstatus_mstatusOld_1_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_tw = next_csr_mstatus_mstatusOld_1_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_38 = next_csr_mstatus_mstatusOld_1_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_tvm = next_csr_mstatus_mstatusOld_1_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_37 = next_csr_mstatus_mstatusOld_1_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_hi_lo_hi_1 = {next_csr_mstatus_mstatusOld_1_tw,
    next_csr_mstatus_mstatusOld_1_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_mxr = next_csr_mstatus_mstatusOld_1_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_36 = next_csr_mstatus_mstatusOld_1_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_hi_hi_lo_1 = {next_csr_mstatus_mstatusOld_1_tw,
    next_csr_mstatus_mstatusOld_1_tvm,next_csr_mstatus_mstatusOld_1_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_sd = next_csr_mstatus_mstatusOld_1_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_41 = next_csr_mstatus_mstatusOld_1_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_WIRE_2_pad0 = next_csr_mstatus_mstatusOld_1_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_T_40 = next_csr_mstatus_mstatusOld_1_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusNew_hi_hi_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_sd,
    next_csr_mstatus_mstatusOld_1_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_2_tsr = next_csr_mstatus_mstatusOld_1_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_39 = next_csr_mstatus_mstatusOld_1_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [9:0] next_csr_mstatus_mstatusNew_hi_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_sd,
    next_csr_mstatus_mstatusOld_1_pad0,next_csr_mstatus_mstatusOld_1_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [12:0] next_csr_mstatus_mstatusNew_hi_hi_1 = {next_csr_mstatus_mstatusOld_1_sd,next_csr_mstatus_mstatusOld_1_pad0
    ,next_csr_mstatus_mstatusOld_1_tsr,next_csr_mstatus_mstatusOld_1_tw,next_csr_mstatus_mstatusOld_1_tvm,
    next_csr_mstatus_mstatusOld_1_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [20:0] next_csr_mstatus_mstatusNew_hi_1 = {next_csr_mstatus_mstatusOld_1_sd,next_csr_mstatus_mstatusOld_1_pad0,
    next_csr_mstatus_mstatusOld_1_tsr,next_csr_mstatus_mstatusOld_1_tw,next_csr_mstatus_mstatusOld_1_tvm,
    next_csr_mstatus_mstatusOld_1_mxr,next_csr_mstatus_mstatusNew_hi_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [31:0] _next_csr_mstatus_mstatusNew_T_4 = {next_csr_mstatus_mstatusOld_1_sd,next_csr_mstatus_mstatusOld_1_pad0,
    next_csr_mstatus_mstatusOld_1_tsr,next_csr_mstatus_mstatusOld_1_tw,next_csr_mstatus_mstatusOld_1_tvm,
    next_csr_mstatus_mstatusOld_1_mxr,next_csr_mstatus_mstatusNew_hi_lo_1,next_csr_mstatus_mstatusNew_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [30:0] _next_csr_mstatus_mstatusNew_T_5 = _next_csr_mstatus_mstatusNew_T_4[30:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:72]
  wire [31:0] next_csr_mstatus_mstatusNew_1 = {next_csr_mstatus_mstatusOld_1_fs == 2'h3,_next_csr_mstatus_mstatusNew_T_4
    [30:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [31:0] _GEN_5191 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_1 : _GEN_5139; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_951 = csrAddr == 12'h340; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_952 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mscratch_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mscratch_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mscratch_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5192 = csrAddr == 12'h340 ? _T_942 : _GEN_5140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_953 = csrAddr == 12'h305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_954 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtvec_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtvec_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mtvec_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5193 = csrAddr == 12'h305 ? _T_942 : _GEN_5141; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_955 = csrAddr == 12'h306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_956 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcounteren_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcounteren_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mcounteren_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5194 = csrAddr == 12'h306 ? _T_942 : _GEN_5142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_957 = csrAddr == 12'h344; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [10:0] _next_csr_mip_T_4 = 11'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mip_T_5 = io_now_csr_mip & 32'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mip_T_6 = _T_942 & 32'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [31:0] _next_csr_mip_T_7 = _next_csr_mip_T_1 | _next_csr_mip_T_6; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [31:0] _GEN_5195 = csrAddr == 12'h344 ? _next_csr_mip_T_7 : _GEN_5143; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_958 = csrAddr == 12'h304; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_959 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mie_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mie_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mie_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5196 = csrAddr == 12'h304 ? _T_942 : _GEN_5144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _T_961 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire  _T_962 = csrAddr == 12'h342; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_963 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_6 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_7 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcause_T_8 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcause_T_9 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_10 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mcause_T_11 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5198 = csrAddr == 12'h342 ? _T_942 : _GEN_5146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_964 = csrAddr == 12'h343; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_965 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtval_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtval_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_28 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _next_csr_mtval_T_29 = rData_3 | _GEN_31; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [31:0] _GEN_5199 = csrAddr == 12'h343 ? _T_942 : _GEN_5147; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5200 = has_15 ? _GEN_5190 : _GEN_5138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5201 = has_15 ? _GEN_5191 : _GEN_5139; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5202 = has_15 ? _GEN_5192 : _GEN_5140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5203 = has_15 ? _GEN_5193 : _GEN_5141; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5204 = has_15 ? _GEN_5194 : _GEN_5142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5205 = has_15 ? _GEN_5195 : _GEN_5143; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5206 = has_15 ? _GEN_5196 : _GEN_5144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5208 = has_15 ? _GEN_5198 : _GEN_5146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5209 = has_15 ? _GEN_5199 : _GEN_5147; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5212 = _T_1090 ? _GEN_5200 : _GEN_5138; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5213 = _T_1090 ? _GEN_5201 : _GEN_5139; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5214 = _T_1090 ? _GEN_5202 : _GEN_5140; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5215 = _T_1090 ? _GEN_5203 : _GEN_5141; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5216 = _T_1090 ? _GEN_5204 : _GEN_5142; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5217 = _T_1090 ? _GEN_5205 : _GEN_5143; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5218 = _T_1090 ? _GEN_5206 : _GEN_5144; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5220 = _T_1090 ? _GEN_5208 : _GEN_5146; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5221 = _T_1090 ? _GEN_5209 : _GEN_5147; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [31:0] _GEN_5224 = _T_1049 ? _GEN_5154 : _GEN_5106; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5225 = _T_1049 ? _GEN_5155 : _GEN_5107; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5226 = _T_1049 ? _GEN_5156 : _GEN_5108; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5227 = _T_1049 ? _GEN_5157 : _GEN_5109; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5228 = _T_1049 ? _GEN_5158 : _GEN_5110; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5229 = _T_1049 ? _GEN_5159 : _GEN_5111; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5230 = _T_1049 ? _GEN_5160 : _GEN_5112; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5231 = _T_1049 ? _GEN_5161 : _GEN_5113; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5232 = _T_1049 ? _GEN_5162 : _GEN_5114; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5233 = _T_1049 ? _GEN_5163 : _GEN_5115; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5234 = _T_1049 ? _GEN_5164 : _GEN_5116; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5235 = _T_1049 ? _GEN_5165 : _GEN_5117; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5236 = _T_1049 ? _GEN_5166 : _GEN_5118; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5237 = _T_1049 ? _GEN_5167 : _GEN_5119; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5238 = _T_1049 ? _GEN_5168 : _GEN_5120; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5239 = _T_1049 ? _GEN_5169 : _GEN_5121; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5240 = _T_1049 ? _GEN_5170 : _GEN_5122; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5241 = _T_1049 ? _GEN_5171 : _GEN_5123; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5242 = _T_1049 ? _GEN_5172 : _GEN_5124; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5243 = _T_1049 ? _GEN_5173 : _GEN_5125; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5244 = _T_1049 ? _GEN_5174 : _GEN_5126; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5245 = _T_1049 ? _GEN_5175 : _GEN_5127; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5246 = _T_1049 ? _GEN_5176 : _GEN_5128; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5247 = _T_1049 ? _GEN_5177 : _GEN_5129; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5248 = _T_1049 ? _GEN_5178 : _GEN_5130; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5249 = _T_1049 ? _GEN_5179 : _GEN_5131; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5250 = _T_1049 ? _GEN_5180 : _GEN_5132; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5251 = _T_1049 ? _GEN_5181 : _GEN_5133; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5252 = _T_1049 ? _GEN_5182 : _GEN_5134; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5253 = _T_1049 ? _GEN_5183 : _GEN_5135; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5254 = _T_1049 ? _GEN_5184 : _GEN_5136; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5255 = _T_1049 ? _GEN_5185 : _GEN_5137; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5256 = _T_1049 ? _GEN_5212 : _GEN_5138; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5257 = _T_1049 ? _GEN_5213 : _GEN_5139; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5258 = _T_1049 ? _GEN_5214 : _GEN_5140; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5259 = _T_1049 ? _GEN_5215 : _GEN_5141; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5260 = _T_1049 ? _GEN_5216 : _GEN_5142; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5261 = _T_1049 ? _GEN_5217 : _GEN_5143; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5262 = _T_1049 ? _GEN_5218 : _GEN_5144; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5264 = _T_1049 ? _GEN_5220 : _GEN_5146; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [31:0] _GEN_5265 = _T_1049 ? _GEN_5221 : _GEN_5147; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [2:0] _GEN_5271 = _T_927 ? inst[14:12] : _GEN_5099; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5273 = _T_927 ? inst[6:0] : _GEN_5101; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_5278 = _T_927 ? _GEN_5224 : _GEN_5106; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5279 = _T_927 ? _GEN_5225 : _GEN_5107; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5280 = _T_927 ? _GEN_5226 : _GEN_5108; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5281 = _T_927 ? _GEN_5227 : _GEN_5109; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5282 = _T_927 ? _GEN_5228 : _GEN_5110; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5283 = _T_927 ? _GEN_5229 : _GEN_5111; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5284 = _T_927 ? _GEN_5230 : _GEN_5112; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5285 = _T_927 ? _GEN_5231 : _GEN_5113; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5286 = _T_927 ? _GEN_5232 : _GEN_5114; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5287 = _T_927 ? _GEN_5233 : _GEN_5115; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5288 = _T_927 ? _GEN_5234 : _GEN_5116; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5289 = _T_927 ? _GEN_5235 : _GEN_5117; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5290 = _T_927 ? _GEN_5236 : _GEN_5118; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5291 = _T_927 ? _GEN_5237 : _GEN_5119; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5292 = _T_927 ? _GEN_5238 : _GEN_5120; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5293 = _T_927 ? _GEN_5239 : _GEN_5121; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5294 = _T_927 ? _GEN_5240 : _GEN_5122; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5295 = _T_927 ? _GEN_5241 : _GEN_5123; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5296 = _T_927 ? _GEN_5242 : _GEN_5124; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5297 = _T_927 ? _GEN_5243 : _GEN_5125; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5298 = _T_927 ? _GEN_5244 : _GEN_5126; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5299 = _T_927 ? _GEN_5245 : _GEN_5127; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5300 = _T_927 ? _GEN_5246 : _GEN_5128; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5301 = _T_927 ? _GEN_5247 : _GEN_5129; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5302 = _T_927 ? _GEN_5248 : _GEN_5130; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5303 = _T_927 ? _GEN_5249 : _GEN_5131; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5304 = _T_927 ? _GEN_5250 : _GEN_5132; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5305 = _T_927 ? _GEN_5251 : _GEN_5133; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5306 = _T_927 ? _GEN_5252 : _GEN_5134; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5307 = _T_927 ? _GEN_5253 : _GEN_5135; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5308 = _T_927 ? _GEN_5254 : _GEN_5136; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5309 = _T_927 ? _GEN_5255 : _GEN_5137; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5310 = _T_927 ? _GEN_5256 : _GEN_5138; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5311 = _T_927 ? _GEN_5257 : _GEN_5139; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5312 = _T_927 ? _GEN_5258 : _GEN_5140; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5313 = _T_927 ? _GEN_5259 : _GEN_5141; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5314 = _T_927 ? _GEN_5260 : _GEN_5142; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5315 = _T_927 ? _GEN_5261 : _GEN_5143; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5316 = _T_927 ? _GEN_5262 : _GEN_5144; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5318 = _T_927 ? _GEN_5264 : _GEN_5146; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [31:0] _GEN_5319 = _T_927 ? _GEN_5265 : _GEN_5147; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [2:0] _funct3_T_69 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_971 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _next_reg_has_T_54 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_55 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_56 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_57 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_58 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_59 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_60 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_61 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_62 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_63 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_64 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_65 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_66 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_67 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_68 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_69 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_70 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_71 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_72 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_73 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_74 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_75 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_76 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_77 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_78 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_79 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_80 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  next_reg_has_2 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_nowCSR_T_54 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_55 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_56 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_57 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_58 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_59 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_60 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_61 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_62 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_63 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_64 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_65 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_66 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_67 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_68 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_69 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_70 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_71 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_72 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_73 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_74 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_75 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_76 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_77 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_78 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_79 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_80 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] next_reg_nowCSR_2 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rmask_T_82 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_83 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_84 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_85 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_86 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_87 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_88 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_89 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_90 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_91 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_92 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_93 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_94 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_95 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _next_reg_rmask_T_96 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_97 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_98 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_99 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_100 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_101 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_102 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_103 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_104 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_105 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_106 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_107 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_108 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_109 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_110 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_111 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_112 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_113 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_114 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_115 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_116 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_117 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_118 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_119 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_120 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_121 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_122 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] next_reg_rmask_2 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_T_191 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] _next_reg_rData_T_12 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rData_T_13 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5322 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire  _next_reg_T_192 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_193 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _next_reg_rData_T_14 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _next_reg_rData_T_15 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _next_reg_rData_T_16 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _next_reg_rData_T_17 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [31:0] _GEN_5323 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5324 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_194 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] next_reg_rData_2 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5325 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_T_195 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_rd_44 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5326 = 5'h0 == rd ? rData_3 : _GEN_5278; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5327 = 5'h1 == rd ? rData_3 : _GEN_5279; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5328 = 5'h2 == rd ? rData_3 : _GEN_5280; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5329 = 5'h3 == rd ? rData_3 : _GEN_5281; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5330 = 5'h4 == rd ? rData_3 : _GEN_5282; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5331 = 5'h5 == rd ? rData_3 : _GEN_5283; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5332 = 5'h6 == rd ? rData_3 : _GEN_5284; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5333 = 5'h7 == rd ? rData_3 : _GEN_5285; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5334 = 5'h8 == rd ? rData_3 : _GEN_5286; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5335 = 5'h9 == rd ? rData_3 : _GEN_5287; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5336 = 5'ha == rd ? rData_3 : _GEN_5288; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5337 = 5'hb == rd ? rData_3 : _GEN_5289; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5338 = 5'hc == rd ? rData_3 : _GEN_5290; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5339 = 5'hd == rd ? rData_3 : _GEN_5291; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5340 = 5'he == rd ? rData_3 : _GEN_5292; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5341 = 5'hf == rd ? rData_3 : _GEN_5293; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5342 = 5'h10 == rd ? rData_3 : _GEN_5294; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5343 = 5'h11 == rd ? rData_3 : _GEN_5295; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5344 = 5'h12 == rd ? rData_3 : _GEN_5296; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5345 = 5'h13 == rd ? rData_3 : _GEN_5297; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5346 = 5'h14 == rd ? rData_3 : _GEN_5298; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5347 = 5'h15 == rd ? rData_3 : _GEN_5299; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5348 = 5'h16 == rd ? rData_3 : _GEN_5300; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5349 = 5'h17 == rd ? rData_3 : _GEN_5301; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5350 = 5'h18 == rd ? rData_3 : _GEN_5302; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5351 = 5'h19 == rd ? rData_3 : _GEN_5303; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5352 = 5'h1a == rd ? rData_3 : _GEN_5304; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5353 = 5'h1b == rd ? rData_3 : _GEN_5305; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5354 = 5'h1c == rd ? rData_3 : _GEN_5306; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5355 = 5'h1d == rd ? rData_3 : _GEN_5307; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5356 = 5'h1e == rd ? rData_3 : _GEN_5308; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [31:0] _GEN_5357 = 5'h1f == rd ? rData_3 : _GEN_5309; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire  _T_979 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_983 = csrAddr == 12'h301; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_984 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_misa_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_misa_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_misa_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5362 = csrAddr == 12'h301 ? _T_982 : _GEN_5310; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_985 = csrAddr == 12'hf11; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_986 = csrAddr == 12'hf12; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_987 = csrAddr == 12'hf13; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_988 = csrAddr == 12'hf14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_989 = csrAddr == 12'h300; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_990 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_14 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_15 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mstatus_T_16 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mstatus_T_17 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_18 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mstatus_T_19 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mstatus_mstatusOld_WIRE_5 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire  next_csr_mstatus_mstatusOld_2_pad4 = _T_982[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sie = _T_982[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_pad3 = _T_982[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mie = _T_982[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_pad2 = _T_982[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_spie = _T_982[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_ube = _T_982[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mpie = _T_982[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_spp = _T_982[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_vs = _T_982[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_mpp = _T_982[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_fs = _T_982[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_xs = _T_982[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mprv = _T_982[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sum = _T_982[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mxr = _T_982[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_tvm = _T_982[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_tw = _T_982[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_tsr = _T_982[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] next_csr_mstatus_mstatusOld_2_pad0 = _T_982[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sd = _T_982[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_4_fs = next_csr_mstatus_mstatusOld_2_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_53 = next_csr_mstatus_mstatusOld_2_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusNew_T_6 = next_csr_mstatus_mstatusOld_2_fs == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:42]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_sie = next_csr_mstatus_mstatusOld_2_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_43 = next_csr_mstatus_mstatusOld_2_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_pad4 = next_csr_mstatus_mstatusOld_2_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_42 = next_csr_mstatus_mstatusOld_2_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_lo_2 = {next_csr_mstatus_mstatusOld_2_sie,
    next_csr_mstatus_mstatusOld_2_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_pad2 = next_csr_mstatus_mstatusOld_2_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_46 = next_csr_mstatus_mstatusOld_2_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_mie = next_csr_mstatus_mstatusOld_2_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_45 = next_csr_mstatus_mstatusOld_2_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_pad2,
    next_csr_mstatus_mstatusOld_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_pad3 = next_csr_mstatus_mstatusOld_2_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_44 = next_csr_mstatus_mstatusOld_2_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_lo_hi_2 = {next_csr_mstatus_mstatusOld_2_pad2,
    next_csr_mstatus_mstatusOld_2_mie,next_csr_mstatus_mstatusOld_2_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [4:0] next_csr_mstatus_mstatusNew_lo_lo_2 = {next_csr_mstatus_mstatusOld_2_pad2,next_csr_mstatus_mstatusOld_2_mie
    ,next_csr_mstatus_mstatusOld_2_pad3,next_csr_mstatus_mstatusOld_2_sie,next_csr_mstatus_mstatusOld_2_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_ube = next_csr_mstatus_mstatusOld_2_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_48 = next_csr_mstatus_mstatusOld_2_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_spie = next_csr_mstatus_mstatusOld_2_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_47 = next_csr_mstatus_mstatusOld_2_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_hi_lo_2 = {next_csr_mstatus_mstatusOld_2_ube,
    next_csr_mstatus_mstatusOld_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_4_vs = next_csr_mstatus_mstatusOld_2_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_51 = next_csr_mstatus_mstatusOld_2_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_spp = next_csr_mstatus_mstatusOld_2_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_50 = next_csr_mstatus_mstatusOld_2_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_hi_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_vs,
    next_csr_mstatus_mstatusOld_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_mpie = next_csr_mstatus_mstatusOld_2_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_49 = next_csr_mstatus_mstatusOld_2_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_lo_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_vs,
    next_csr_mstatus_mstatusOld_2_spp,next_csr_mstatus_mstatusOld_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_hi_2 = {next_csr_mstatus_mstatusOld_2_vs,next_csr_mstatus_mstatusOld_2_spp,
    next_csr_mstatus_mstatusOld_2_mpie,next_csr_mstatus_mstatusOld_2_ube,next_csr_mstatus_mstatusOld_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [10:0] next_csr_mstatus_mstatusNew_lo_2 = {next_csr_mstatus_mstatusOld_2_vs,next_csr_mstatus_mstatusOld_2_spp,
    next_csr_mstatus_mstatusOld_2_mpie,next_csr_mstatus_mstatusOld_2_ube,next_csr_mstatus_mstatusOld_2_spie,
    next_csr_mstatus_mstatusOld_2_pad2,next_csr_mstatus_mstatusOld_2_mie,next_csr_mstatus_mstatusOld_2_pad3,
    next_csr_mstatus_mstatusOld_2_sie,next_csr_mstatus_mstatusOld_2_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_4_mpp = next_csr_mstatus_mstatusOld_2_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_52 = next_csr_mstatus_mstatusOld_2_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_lo_2 = {next_csr_mstatus_mstatusOld_2_fs,
    next_csr_mstatus_mstatusOld_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_sum = next_csr_mstatus_mstatusOld_2_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_56 = next_csr_mstatus_mstatusOld_2_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_mprv = next_csr_mstatus_mstatusOld_2_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_55 = next_csr_mstatus_mstatusOld_2_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_lo_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_sum,
    next_csr_mstatus_mstatusOld_2_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_4_xs = next_csr_mstatus_mstatusOld_2_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_54 = next_csr_mstatus_mstatusOld_2_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_hi_2 = {next_csr_mstatus_mstatusOld_2_sum,
    next_csr_mstatus_mstatusOld_2_mprv,next_csr_mstatus_mstatusOld_2_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [7:0] next_csr_mstatus_mstatusNew_hi_lo_2 = {next_csr_mstatus_mstatusOld_2_sum,next_csr_mstatus_mstatusOld_2_mprv
    ,next_csr_mstatus_mstatusOld_2_xs,next_csr_mstatus_mstatusOld_2_fs,next_csr_mstatus_mstatusOld_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_tw = next_csr_mstatus_mstatusOld_2_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_59 = next_csr_mstatus_mstatusOld_2_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_tvm = next_csr_mstatus_mstatusOld_2_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_58 = next_csr_mstatus_mstatusOld_2_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_hi_lo_hi_2 = {next_csr_mstatus_mstatusOld_2_tw,
    next_csr_mstatus_mstatusOld_2_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_mxr = next_csr_mstatus_mstatusOld_2_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_57 = next_csr_mstatus_mstatusOld_2_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_hi_hi_lo_2 = {next_csr_mstatus_mstatusOld_2_tw,
    next_csr_mstatus_mstatusOld_2_tvm,next_csr_mstatus_mstatusOld_2_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_sd = next_csr_mstatus_mstatusOld_2_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_62 = next_csr_mstatus_mstatusOld_2_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_WIRE_4_pad0 = next_csr_mstatus_mstatusOld_2_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_T_61 = next_csr_mstatus_mstatusOld_2_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusNew_hi_hi_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_sd,
    next_csr_mstatus_mstatusOld_2_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_4_tsr = next_csr_mstatus_mstatusOld_2_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_60 = next_csr_mstatus_mstatusOld_2_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [9:0] next_csr_mstatus_mstatusNew_hi_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_sd,
    next_csr_mstatus_mstatusOld_2_pad0,next_csr_mstatus_mstatusOld_2_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [12:0] next_csr_mstatus_mstatusNew_hi_hi_2 = {next_csr_mstatus_mstatusOld_2_sd,next_csr_mstatus_mstatusOld_2_pad0
    ,next_csr_mstatus_mstatusOld_2_tsr,next_csr_mstatus_mstatusOld_2_tw,next_csr_mstatus_mstatusOld_2_tvm,
    next_csr_mstatus_mstatusOld_2_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [20:0] next_csr_mstatus_mstatusNew_hi_2 = {next_csr_mstatus_mstatusOld_2_sd,next_csr_mstatus_mstatusOld_2_pad0,
    next_csr_mstatus_mstatusOld_2_tsr,next_csr_mstatus_mstatusOld_2_tw,next_csr_mstatus_mstatusOld_2_tvm,
    next_csr_mstatus_mstatusOld_2_mxr,next_csr_mstatus_mstatusNew_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [31:0] _next_csr_mstatus_mstatusNew_T_7 = {next_csr_mstatus_mstatusOld_2_sd,next_csr_mstatus_mstatusOld_2_pad0,
    next_csr_mstatus_mstatusOld_2_tsr,next_csr_mstatus_mstatusOld_2_tw,next_csr_mstatus_mstatusOld_2_tvm,
    next_csr_mstatus_mstatusOld_2_mxr,next_csr_mstatus_mstatusNew_hi_lo_2,next_csr_mstatus_mstatusNew_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [30:0] _next_csr_mstatus_mstatusNew_T_8 = _next_csr_mstatus_mstatusNew_T_7[30:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:72]
  wire [31:0] next_csr_mstatus_mstatusNew_2 = {next_csr_mstatus_mstatusOld_2_fs == 2'h3,_next_csr_mstatus_mstatusNew_T_7
    [30:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [31:0] _GEN_5363 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_2 : _GEN_5311; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_991 = csrAddr == 12'h340; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_992 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mscratch_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mscratch_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mscratch_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5364 = csrAddr == 12'h340 ? _T_982 : _GEN_5312; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_993 = csrAddr == 12'h305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_994 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtvec_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtvec_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mtvec_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5365 = csrAddr == 12'h305 ? _T_982 : _GEN_5313; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_995 = csrAddr == 12'h306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_996 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcounteren_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcounteren_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mcounteren_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5366 = csrAddr == 12'h306 ? _T_982 : _GEN_5314; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_997 = csrAddr == 12'h344; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [10:0] _next_csr_mip_T_8 = 11'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mip_T_9 = io_now_csr_mip & 32'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mip_T_10 = _T_982 & 32'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [31:0] _next_csr_mip_T_11 = _next_csr_mip_T_1 | _next_csr_mip_T_10; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [31:0] _GEN_5367 = csrAddr == 12'h344 ? _next_csr_mip_T_11 : _GEN_5315; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_998 = csrAddr == 12'h304; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_999 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mie_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mie_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mie_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5368 = csrAddr == 12'h304 ? _T_982 : _GEN_5316; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _T_1001 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire  _T_1002 = csrAddr == 12'h342; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1003 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_12 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_13 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcause_T_14 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcause_T_15 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_16 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mcause_T_17 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5370 = csrAddr == 12'h342 ? _T_982 : _GEN_5318; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1004 = csrAddr == 12'h343; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1005 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtval_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtval_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_34 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _next_csr_mtval_T_35 = rData_3 & _T_981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [31:0] _GEN_5371 = csrAddr == 12'h343 ? _T_982 : _GEN_5319; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5372 = has_15 ? _GEN_5362 : _GEN_5310; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5373 = has_15 ? _GEN_5363 : _GEN_5311; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5374 = has_15 ? _GEN_5364 : _GEN_5312; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5375 = has_15 ? _GEN_5365 : _GEN_5313; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5376 = has_15 ? _GEN_5366 : _GEN_5314; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5377 = has_15 ? _GEN_5367 : _GEN_5315; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5378 = has_15 ? _GEN_5368 : _GEN_5316; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5380 = has_15 ? _GEN_5370 : _GEN_5318; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5381 = has_15 ? _GEN_5371 : _GEN_5319; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5384 = _T_1090 ? _GEN_5372 : _GEN_5310; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5385 = _T_1090 ? _GEN_5373 : _GEN_5311; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5386 = _T_1090 ? _GEN_5374 : _GEN_5312; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5387 = _T_1090 ? _GEN_5375 : _GEN_5313; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5388 = _T_1090 ? _GEN_5376 : _GEN_5314; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5389 = _T_1090 ? _GEN_5377 : _GEN_5315; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5390 = _T_1090 ? _GEN_5378 : _GEN_5316; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5392 = _T_1090 ? _GEN_5380 : _GEN_5318; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5393 = _T_1090 ? _GEN_5381 : _GEN_5319; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [31:0] _GEN_5396 = _T_1089 ? _GEN_5326 : _GEN_5278; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5397 = _T_1089 ? _GEN_5327 : _GEN_5279; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5398 = _T_1089 ? _GEN_5328 : _GEN_5280; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5399 = _T_1089 ? _GEN_5329 : _GEN_5281; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5400 = _T_1089 ? _GEN_5330 : _GEN_5282; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5401 = _T_1089 ? _GEN_5331 : _GEN_5283; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5402 = _T_1089 ? _GEN_5332 : _GEN_5284; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5403 = _T_1089 ? _GEN_5333 : _GEN_5285; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5404 = _T_1089 ? _GEN_5334 : _GEN_5286; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5405 = _T_1089 ? _GEN_5335 : _GEN_5287; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5406 = _T_1089 ? _GEN_5336 : _GEN_5288; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5407 = _T_1089 ? _GEN_5337 : _GEN_5289; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5408 = _T_1089 ? _GEN_5338 : _GEN_5290; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5409 = _T_1089 ? _GEN_5339 : _GEN_5291; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5410 = _T_1089 ? _GEN_5340 : _GEN_5292; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5411 = _T_1089 ? _GEN_5341 : _GEN_5293; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5412 = _T_1089 ? _GEN_5342 : _GEN_5294; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5413 = _T_1089 ? _GEN_5343 : _GEN_5295; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5414 = _T_1089 ? _GEN_5344 : _GEN_5296; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5415 = _T_1089 ? _GEN_5345 : _GEN_5297; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5416 = _T_1089 ? _GEN_5346 : _GEN_5298; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5417 = _T_1089 ? _GEN_5347 : _GEN_5299; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5418 = _T_1089 ? _GEN_5348 : _GEN_5300; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5419 = _T_1089 ? _GEN_5349 : _GEN_5301; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5420 = _T_1089 ? _GEN_5350 : _GEN_5302; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5421 = _T_1089 ? _GEN_5351 : _GEN_5303; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5422 = _T_1089 ? _GEN_5352 : _GEN_5304; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5423 = _T_1089 ? _GEN_5353 : _GEN_5305; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5424 = _T_1089 ? _GEN_5354 : _GEN_5306; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5425 = _T_1089 ? _GEN_5355 : _GEN_5307; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5426 = _T_1089 ? _GEN_5356 : _GEN_5308; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5427 = _T_1089 ? _GEN_5357 : _GEN_5309; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5428 = _T_1089 ? _GEN_5384 : _GEN_5310; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5429 = _T_1089 ? _GEN_5385 : _GEN_5311; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5430 = _T_1089 ? _GEN_5386 : _GEN_5312; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5431 = _T_1089 ? _GEN_5387 : _GEN_5313; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5432 = _T_1089 ? _GEN_5388 : _GEN_5314; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5433 = _T_1089 ? _GEN_5389 : _GEN_5315; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5434 = _T_1089 ? _GEN_5390 : _GEN_5316; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5436 = _T_1089 ? _GEN_5392 : _GEN_5318; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [31:0] _GEN_5437 = _T_1089 ? _GEN_5393 : _GEN_5319; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [2:0] _GEN_5443 = _T_967 ? inst[14:12] : _GEN_5271; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5445 = _T_967 ? inst[6:0] : _GEN_5273; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_5450 = _T_967 ? _GEN_5396 : _GEN_5278; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5451 = _T_967 ? _GEN_5397 : _GEN_5279; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5452 = _T_967 ? _GEN_5398 : _GEN_5280; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5453 = _T_967 ? _GEN_5399 : _GEN_5281; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5454 = _T_967 ? _GEN_5400 : _GEN_5282; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5455 = _T_967 ? _GEN_5401 : _GEN_5283; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5456 = _T_967 ? _GEN_5402 : _GEN_5284; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5457 = _T_967 ? _GEN_5403 : _GEN_5285; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5458 = _T_967 ? _GEN_5404 : _GEN_5286; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5459 = _T_967 ? _GEN_5405 : _GEN_5287; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5460 = _T_967 ? _GEN_5406 : _GEN_5288; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5461 = _T_967 ? _GEN_5407 : _GEN_5289; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5462 = _T_967 ? _GEN_5408 : _GEN_5290; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5463 = _T_967 ? _GEN_5409 : _GEN_5291; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5464 = _T_967 ? _GEN_5410 : _GEN_5292; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5465 = _T_967 ? _GEN_5411 : _GEN_5293; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5466 = _T_967 ? _GEN_5412 : _GEN_5294; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5467 = _T_967 ? _GEN_5413 : _GEN_5295; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5468 = _T_967 ? _GEN_5414 : _GEN_5296; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5469 = _T_967 ? _GEN_5415 : _GEN_5297; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5470 = _T_967 ? _GEN_5416 : _GEN_5298; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5471 = _T_967 ? _GEN_5417 : _GEN_5299; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5472 = _T_967 ? _GEN_5418 : _GEN_5300; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5473 = _T_967 ? _GEN_5419 : _GEN_5301; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5474 = _T_967 ? _GEN_5420 : _GEN_5302; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5475 = _T_967 ? _GEN_5421 : _GEN_5303; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5476 = _T_967 ? _GEN_5422 : _GEN_5304; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5477 = _T_967 ? _GEN_5423 : _GEN_5305; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5478 = _T_967 ? _GEN_5424 : _GEN_5306; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5479 = _T_967 ? _GEN_5425 : _GEN_5307; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5480 = _T_967 ? _GEN_5426 : _GEN_5308; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5481 = _T_967 ? _GEN_5427 : _GEN_5309; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5482 = _T_967 ? _GEN_5428 : _GEN_5310; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5483 = _T_967 ? _GEN_5429 : _GEN_5311; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5484 = _T_967 ? _GEN_5430 : _GEN_5312; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5485 = _T_967 ? _GEN_5431 : _GEN_5313; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5486 = _T_967 ? _GEN_5432 : _GEN_5314; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5487 = _T_967 ? _GEN_5433 : _GEN_5315; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5488 = _T_967 ? _GEN_5434 : _GEN_5316; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5490 = _T_967 ? _GEN_5436 : _GEN_5318; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [31:0] _GEN_5491 = _T_967 ? _GEN_5437 : _GEN_5319; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [2:0] _funct3_T_70 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_1011 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _T_1015 = rd != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:17]
  wire  _next_reg_has_T_81 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_82 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_83 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_84 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_85 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_86 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_87 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_88 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_89 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_90 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_91 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_92 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_93 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_94 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_95 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_96 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_97 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_98 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_99 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_100 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_101 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_102 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_103 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_104 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_105 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_106 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_107 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  next_reg_has_3 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_nowCSR_T_81 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_82 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_83 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_84 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_85 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_86 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_87 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_88 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_89 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_90 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_91 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_92 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_93 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_94 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_95 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_96 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_97 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_98 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_99 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_100 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_101 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_102 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_103 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_104 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_105 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_106 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_107 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] next_reg_nowCSR_3 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rmask_T_123 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_124 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_125 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_126 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_127 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_128 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_129 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_130 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_131 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_132 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_133 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_134 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_135 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_136 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _next_reg_rmask_T_137 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_138 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_139 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_140 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_141 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_142 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_143 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_144 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_145 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_146 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_147 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_148 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_149 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_150 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_151 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_152 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_153 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_154 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_155 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_156 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_157 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_158 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_159 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_160 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_161 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_162 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_163 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] next_reg_rmask_3 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_T_196 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] _next_reg_rData_T_18 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rData_T_19 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5494 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire  _next_reg_T_197 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_198 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _next_reg_rData_T_20 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _next_reg_rData_T_21 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _next_reg_rData_T_22 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _next_reg_rData_T_23 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [31:0] _GEN_5495 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5496 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_199 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] next_reg_rData_3 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5497 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_T_200 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_rd_45 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5498 = 5'h0 == rd ? rData_3 : _GEN_5450; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5499 = 5'h1 == rd ? rData_3 : _GEN_5451; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5500 = 5'h2 == rd ? rData_3 : _GEN_5452; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5501 = 5'h3 == rd ? rData_3 : _GEN_5453; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5502 = 5'h4 == rd ? rData_3 : _GEN_5454; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5503 = 5'h5 == rd ? rData_3 : _GEN_5455; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5504 = 5'h6 == rd ? rData_3 : _GEN_5456; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5505 = 5'h7 == rd ? rData_3 : _GEN_5457; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5506 = 5'h8 == rd ? rData_3 : _GEN_5458; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5507 = 5'h9 == rd ? rData_3 : _GEN_5459; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5508 = 5'ha == rd ? rData_3 : _GEN_5460; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5509 = 5'hb == rd ? rData_3 : _GEN_5461; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5510 = 5'hc == rd ? rData_3 : _GEN_5462; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5511 = 5'hd == rd ? rData_3 : _GEN_5463; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5512 = 5'he == rd ? rData_3 : _GEN_5464; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5513 = 5'hf == rd ? rData_3 : _GEN_5465; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5514 = 5'h10 == rd ? rData_3 : _GEN_5466; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5515 = 5'h11 == rd ? rData_3 : _GEN_5467; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5516 = 5'h12 == rd ? rData_3 : _GEN_5468; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5517 = 5'h13 == rd ? rData_3 : _GEN_5469; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5518 = 5'h14 == rd ? rData_3 : _GEN_5470; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5519 = 5'h15 == rd ? rData_3 : _GEN_5471; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5520 = 5'h16 == rd ? rData_3 : _GEN_5472; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5521 = 5'h17 == rd ? rData_3 : _GEN_5473; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5522 = 5'h18 == rd ? rData_3 : _GEN_5474; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5523 = 5'h19 == rd ? rData_3 : _GEN_5475; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5524 = 5'h1a == rd ? rData_3 : _GEN_5476; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5525 = 5'h1b == rd ? rData_3 : _GEN_5477; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5526 = 5'h1c == rd ? rData_3 : _GEN_5478; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5527 = 5'h1d == rd ? rData_3 : _GEN_5479; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5528 = 5'h1e == rd ? rData_3 : _GEN_5480; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5529 = 5'h1f == rd ? rData_3 : _GEN_5481; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [31:0] _GEN_5530 = _T_902 ? _GEN_5498 : _GEN_5450; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5531 = _T_902 ? _GEN_5499 : _GEN_5451; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5532 = _T_902 ? _GEN_5500 : _GEN_5452; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5533 = _T_902 ? _GEN_5501 : _GEN_5453; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5534 = _T_902 ? _GEN_5502 : _GEN_5454; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5535 = _T_902 ? _GEN_5503 : _GEN_5455; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5536 = _T_902 ? _GEN_5504 : _GEN_5456; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5537 = _T_902 ? _GEN_5505 : _GEN_5457; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5538 = _T_902 ? _GEN_5506 : _GEN_5458; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5539 = _T_902 ? _GEN_5507 : _GEN_5459; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5540 = _T_902 ? _GEN_5508 : _GEN_5460; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5541 = _T_902 ? _GEN_5509 : _GEN_5461; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5542 = _T_902 ? _GEN_5510 : _GEN_5462; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5543 = _T_902 ? _GEN_5511 : _GEN_5463; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5544 = _T_902 ? _GEN_5512 : _GEN_5464; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5545 = _T_902 ? _GEN_5513 : _GEN_5465; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5546 = _T_902 ? _GEN_5514 : _GEN_5466; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5547 = _T_902 ? _GEN_5515 : _GEN_5467; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5548 = _T_902 ? _GEN_5516 : _GEN_5468; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5549 = _T_902 ? _GEN_5517 : _GEN_5469; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5550 = _T_902 ? _GEN_5518 : _GEN_5470; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5551 = _T_902 ? _GEN_5519 : _GEN_5471; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5552 = _T_902 ? _GEN_5520 : _GEN_5472; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5553 = _T_902 ? _GEN_5521 : _GEN_5473; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5554 = _T_902 ? _GEN_5522 : _GEN_5474; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5555 = _T_902 ? _GEN_5523 : _GEN_5475; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5556 = _T_902 ? _GEN_5524 : _GEN_5476; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5557 = _T_902 ? _GEN_5525 : _GEN_5477; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5558 = _T_902 ? _GEN_5526 : _GEN_5478; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5559 = _T_902 ? _GEN_5527 : _GEN_5479; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5560 = _T_902 ? _GEN_5528 : _GEN_5480; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [31:0] _GEN_5561 = _T_902 ? _GEN_5529 : _GEN_5481; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire  _T_1017 = csrAddr == 12'h301; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1018 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_misa_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_misa_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_misa_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5562 = csrAddr == 12'h301 ? _T_1096 : _GEN_5482; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1019 = csrAddr == 12'hf11; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1020 = csrAddr == 12'hf12; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1021 = csrAddr == 12'hf13; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1022 = csrAddr == 12'hf14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1023 = csrAddr == 12'h300; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1024 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_20 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_21 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mstatus_T_22 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mstatus_T_23 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_24 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mstatus_T_25 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mstatus_mstatusOld_WIRE_7 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  next_csr_mstatus_mstatusOld_3_pad4 = _T_1096[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sie = _T_1096[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_pad3 = _T_1096[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mie = _T_1096[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_pad2 = _T_1096[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_spie = _T_1096[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_ube = _T_1096[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mpie = _T_1096[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_spp = _T_1096[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_vs = _T_1096[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_mpp = _T_1096[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_fs = _T_1096[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_xs = _T_1096[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mprv = _T_1096[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sum = _T_1096[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mxr = _T_1096[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_tvm = _T_1096[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_tw = _T_1096[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_tsr = _T_1096[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] next_csr_mstatus_mstatusOld_3_pad0 = _T_1096[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sd = _T_1096[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_6_fs = next_csr_mstatus_mstatusOld_3_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_74 = next_csr_mstatus_mstatusOld_3_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusNew_T_9 = next_csr_mstatus_mstatusOld_3_fs == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:42]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_sie = next_csr_mstatus_mstatusOld_3_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_64 = next_csr_mstatus_mstatusOld_3_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_pad4 = next_csr_mstatus_mstatusOld_3_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_63 = next_csr_mstatus_mstatusOld_3_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_lo_3 = {next_csr_mstatus_mstatusOld_3_sie,
    next_csr_mstatus_mstatusOld_3_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_pad2 = next_csr_mstatus_mstatusOld_3_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_67 = next_csr_mstatus_mstatusOld_3_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_mie = next_csr_mstatus_mstatusOld_3_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_66 = next_csr_mstatus_mstatusOld_3_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_pad2,
    next_csr_mstatus_mstatusOld_3_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_pad3 = next_csr_mstatus_mstatusOld_3_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_65 = next_csr_mstatus_mstatusOld_3_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_lo_hi_3 = {next_csr_mstatus_mstatusOld_3_pad2,
    next_csr_mstatus_mstatusOld_3_mie,next_csr_mstatus_mstatusOld_3_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [4:0] next_csr_mstatus_mstatusNew_lo_lo_3 = {next_csr_mstatus_mstatusOld_3_pad2,next_csr_mstatus_mstatusOld_3_mie
    ,next_csr_mstatus_mstatusOld_3_pad3,next_csr_mstatus_mstatusOld_3_sie,next_csr_mstatus_mstatusOld_3_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_ube = next_csr_mstatus_mstatusOld_3_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_69 = next_csr_mstatus_mstatusOld_3_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_spie = next_csr_mstatus_mstatusOld_3_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_68 = next_csr_mstatus_mstatusOld_3_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_hi_lo_3 = {next_csr_mstatus_mstatusOld_3_ube,
    next_csr_mstatus_mstatusOld_3_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_6_vs = next_csr_mstatus_mstatusOld_3_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_72 = next_csr_mstatus_mstatusOld_3_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_spp = next_csr_mstatus_mstatusOld_3_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_71 = next_csr_mstatus_mstatusOld_3_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_hi_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_vs,
    next_csr_mstatus_mstatusOld_3_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_mpie = next_csr_mstatus_mstatusOld_3_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_70 = next_csr_mstatus_mstatusOld_3_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_lo_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_vs,
    next_csr_mstatus_mstatusOld_3_spp,next_csr_mstatus_mstatusOld_3_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_hi_3 = {next_csr_mstatus_mstatusOld_3_vs,next_csr_mstatus_mstatusOld_3_spp,
    next_csr_mstatus_mstatusOld_3_mpie,next_csr_mstatus_mstatusOld_3_ube,next_csr_mstatus_mstatusOld_3_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [10:0] next_csr_mstatus_mstatusNew_lo_3 = {next_csr_mstatus_mstatusOld_3_vs,next_csr_mstatus_mstatusOld_3_spp,
    next_csr_mstatus_mstatusOld_3_mpie,next_csr_mstatus_mstatusOld_3_ube,next_csr_mstatus_mstatusOld_3_spie,
    next_csr_mstatus_mstatusOld_3_pad2,next_csr_mstatus_mstatusOld_3_mie,next_csr_mstatus_mstatusOld_3_pad3,
    next_csr_mstatus_mstatusOld_3_sie,next_csr_mstatus_mstatusOld_3_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_6_mpp = next_csr_mstatus_mstatusOld_3_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_73 = next_csr_mstatus_mstatusOld_3_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_lo_3 = {next_csr_mstatus_mstatusOld_3_fs,
    next_csr_mstatus_mstatusOld_3_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_sum = next_csr_mstatus_mstatusOld_3_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_77 = next_csr_mstatus_mstatusOld_3_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_mprv = next_csr_mstatus_mstatusOld_3_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_76 = next_csr_mstatus_mstatusOld_3_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_lo_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_sum,
    next_csr_mstatus_mstatusOld_3_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_6_xs = next_csr_mstatus_mstatusOld_3_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_75 = next_csr_mstatus_mstatusOld_3_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_hi_3 = {next_csr_mstatus_mstatusOld_3_sum,
    next_csr_mstatus_mstatusOld_3_mprv,next_csr_mstatus_mstatusOld_3_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [7:0] next_csr_mstatus_mstatusNew_hi_lo_3 = {next_csr_mstatus_mstatusOld_3_sum,next_csr_mstatus_mstatusOld_3_mprv
    ,next_csr_mstatus_mstatusOld_3_xs,next_csr_mstatus_mstatusOld_3_fs,next_csr_mstatus_mstatusOld_3_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_tw = next_csr_mstatus_mstatusOld_3_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_80 = next_csr_mstatus_mstatusOld_3_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_tvm = next_csr_mstatus_mstatusOld_3_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_79 = next_csr_mstatus_mstatusOld_3_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_hi_lo_hi_3 = {next_csr_mstatus_mstatusOld_3_tw,
    next_csr_mstatus_mstatusOld_3_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_mxr = next_csr_mstatus_mstatusOld_3_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_78 = next_csr_mstatus_mstatusOld_3_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_hi_hi_lo_3 = {next_csr_mstatus_mstatusOld_3_tw,
    next_csr_mstatus_mstatusOld_3_tvm,next_csr_mstatus_mstatusOld_3_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_sd = next_csr_mstatus_mstatusOld_3_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_83 = next_csr_mstatus_mstatusOld_3_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_WIRE_6_pad0 = next_csr_mstatus_mstatusOld_3_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_T_82 = next_csr_mstatus_mstatusOld_3_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusNew_hi_hi_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_sd,
    next_csr_mstatus_mstatusOld_3_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_6_tsr = next_csr_mstatus_mstatusOld_3_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_81 = next_csr_mstatus_mstatusOld_3_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [9:0] next_csr_mstatus_mstatusNew_hi_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_sd,
    next_csr_mstatus_mstatusOld_3_pad0,next_csr_mstatus_mstatusOld_3_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [12:0] next_csr_mstatus_mstatusNew_hi_hi_3 = {next_csr_mstatus_mstatusOld_3_sd,next_csr_mstatus_mstatusOld_3_pad0
    ,next_csr_mstatus_mstatusOld_3_tsr,next_csr_mstatus_mstatusOld_3_tw,next_csr_mstatus_mstatusOld_3_tvm,
    next_csr_mstatus_mstatusOld_3_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [20:0] next_csr_mstatus_mstatusNew_hi_3 = {next_csr_mstatus_mstatusOld_3_sd,next_csr_mstatus_mstatusOld_3_pad0,
    next_csr_mstatus_mstatusOld_3_tsr,next_csr_mstatus_mstatusOld_3_tw,next_csr_mstatus_mstatusOld_3_tvm,
    next_csr_mstatus_mstatusOld_3_mxr,next_csr_mstatus_mstatusNew_hi_lo_3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [31:0] _next_csr_mstatus_mstatusNew_T_10 = {next_csr_mstatus_mstatusOld_3_sd,next_csr_mstatus_mstatusOld_3_pad0,
    next_csr_mstatus_mstatusOld_3_tsr,next_csr_mstatus_mstatusOld_3_tw,next_csr_mstatus_mstatusOld_3_tvm,
    next_csr_mstatus_mstatusOld_3_mxr,next_csr_mstatus_mstatusNew_hi_lo_3,next_csr_mstatus_mstatusNew_lo_3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [30:0] _next_csr_mstatus_mstatusNew_T_11 = _next_csr_mstatus_mstatusNew_T_10[30:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:72]
  wire [31:0] next_csr_mstatus_mstatusNew_3 = {next_csr_mstatus_mstatusOld_3_fs == 2'h3,
    _next_csr_mstatus_mstatusNew_T_10[30:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [31:0] _GEN_5563 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_3 : _GEN_5483; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1025 = csrAddr == 12'h340; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1026 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mscratch_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mscratch_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mscratch_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5564 = csrAddr == 12'h340 ? _T_1096 : _GEN_5484; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1027 = csrAddr == 12'h305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1028 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtvec_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtvec_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mtvec_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5565 = csrAddr == 12'h305 ? _T_1096 : _GEN_5485; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1029 = csrAddr == 12'h306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1030 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcounteren_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcounteren_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mcounteren_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5566 = csrAddr == 12'h306 ? _T_1096 : _GEN_5486; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1031 = csrAddr == 12'h344; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [10:0] _next_csr_mip_T_12 = 11'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mip_T_13 = io_now_csr_mip & 32'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mip_T_14 = _T_1096 & 32'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [31:0] _next_csr_mip_T_15 = _next_csr_mip_T_1 | _next_csr_mip_T_14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [31:0] _GEN_5567 = csrAddr == 12'h344 ? _next_csr_mip_T_15 : _GEN_5487; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1032 = csrAddr == 12'h304; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1033 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mie_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mie_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mie_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5568 = csrAddr == 12'h304 ? _T_1096 : _GEN_5488; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _T_1035 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire  _T_1036 = csrAddr == 12'h342; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1037 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_18 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_19 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcause_T_20 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcause_T_21 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_22 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mcause_T_23 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5570 = csrAddr == 12'h342 ? _T_1096 : _GEN_5490; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1038 = csrAddr == 12'h343; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1039 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_36 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_37 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtval_T_38 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtval_T_39 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_40 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mtval_T_41 = {27'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_5571 = csrAddr == 12'h343 ? _T_1096 : _GEN_5491; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5572 = has_15 ? _GEN_5562 : _GEN_5482; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5573 = has_15 ? _GEN_5563 : _GEN_5483; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5574 = has_15 ? _GEN_5564 : _GEN_5484; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5575 = has_15 ? _GEN_5565 : _GEN_5485; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5576 = has_15 ? _GEN_5566 : _GEN_5486; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5577 = has_15 ? _GEN_5567 : _GEN_5487; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5578 = has_15 ? _GEN_5568 : _GEN_5488; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5580 = has_15 ? _GEN_5570 : _GEN_5490; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5581 = has_15 ? _GEN_5571 : _GEN_5491; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5584 = _T_1089 ? _GEN_5530 : _GEN_5450; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5585 = _T_1089 ? _GEN_5531 : _GEN_5451; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5586 = _T_1089 ? _GEN_5532 : _GEN_5452; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5587 = _T_1089 ? _GEN_5533 : _GEN_5453; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5588 = _T_1089 ? _GEN_5534 : _GEN_5454; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5589 = _T_1089 ? _GEN_5535 : _GEN_5455; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5590 = _T_1089 ? _GEN_5536 : _GEN_5456; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5591 = _T_1089 ? _GEN_5537 : _GEN_5457; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5592 = _T_1089 ? _GEN_5538 : _GEN_5458; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5593 = _T_1089 ? _GEN_5539 : _GEN_5459; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5594 = _T_1089 ? _GEN_5540 : _GEN_5460; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5595 = _T_1089 ? _GEN_5541 : _GEN_5461; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5596 = _T_1089 ? _GEN_5542 : _GEN_5462; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5597 = _T_1089 ? _GEN_5543 : _GEN_5463; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5598 = _T_1089 ? _GEN_5544 : _GEN_5464; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5599 = _T_1089 ? _GEN_5545 : _GEN_5465; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5600 = _T_1089 ? _GEN_5546 : _GEN_5466; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5601 = _T_1089 ? _GEN_5547 : _GEN_5467; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5602 = _T_1089 ? _GEN_5548 : _GEN_5468; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5603 = _T_1089 ? _GEN_5549 : _GEN_5469; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5604 = _T_1089 ? _GEN_5550 : _GEN_5470; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5605 = _T_1089 ? _GEN_5551 : _GEN_5471; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5606 = _T_1089 ? _GEN_5552 : _GEN_5472; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5607 = _T_1089 ? _GEN_5553 : _GEN_5473; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5608 = _T_1089 ? _GEN_5554 : _GEN_5474; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5609 = _T_1089 ? _GEN_5555 : _GEN_5475; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5610 = _T_1089 ? _GEN_5556 : _GEN_5476; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5611 = _T_1089 ? _GEN_5557 : _GEN_5477; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5612 = _T_1089 ? _GEN_5558 : _GEN_5478; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5613 = _T_1089 ? _GEN_5559 : _GEN_5479; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5614 = _T_1089 ? _GEN_5560 : _GEN_5480; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5615 = _T_1089 ? _GEN_5561 : _GEN_5481; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5616 = _T_1089 ? _GEN_5572 : _GEN_5482; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5617 = _T_1089 ? _GEN_5573 : _GEN_5483; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5618 = _T_1089 ? _GEN_5574 : _GEN_5484; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5619 = _T_1089 ? _GEN_5575 : _GEN_5485; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5620 = _T_1089 ? _GEN_5576 : _GEN_5486; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5621 = _T_1089 ? _GEN_5577 : _GEN_5487; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5622 = _T_1089 ? _GEN_5578 : _GEN_5488; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5624 = _T_1089 ? _GEN_5580 : _GEN_5490; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [31:0] _GEN_5625 = _T_1089 ? _GEN_5581 : _GEN_5491; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [2:0] _GEN_5631 = _T_1007 ? inst[14:12] : _GEN_5443; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5633 = _T_1007 ? inst[6:0] : _GEN_5445; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_5638 = _T_1007 ? _GEN_5584 : _GEN_5450; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5639 = _T_1007 ? _GEN_5585 : _GEN_5451; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5640 = _T_1007 ? _GEN_5586 : _GEN_5452; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5641 = _T_1007 ? _GEN_5587 : _GEN_5453; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5642 = _T_1007 ? _GEN_5588 : _GEN_5454; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5643 = _T_1007 ? _GEN_5589 : _GEN_5455; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5644 = _T_1007 ? _GEN_5590 : _GEN_5456; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5645 = _T_1007 ? _GEN_5591 : _GEN_5457; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5646 = _T_1007 ? _GEN_5592 : _GEN_5458; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5647 = _T_1007 ? _GEN_5593 : _GEN_5459; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5648 = _T_1007 ? _GEN_5594 : _GEN_5460; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5649 = _T_1007 ? _GEN_5595 : _GEN_5461; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5650 = _T_1007 ? _GEN_5596 : _GEN_5462; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5651 = _T_1007 ? _GEN_5597 : _GEN_5463; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5652 = _T_1007 ? _GEN_5598 : _GEN_5464; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5653 = _T_1007 ? _GEN_5599 : _GEN_5465; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5654 = _T_1007 ? _GEN_5600 : _GEN_5466; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5655 = _T_1007 ? _GEN_5601 : _GEN_5467; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5656 = _T_1007 ? _GEN_5602 : _GEN_5468; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5657 = _T_1007 ? _GEN_5603 : _GEN_5469; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5658 = _T_1007 ? _GEN_5604 : _GEN_5470; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5659 = _T_1007 ? _GEN_5605 : _GEN_5471; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5660 = _T_1007 ? _GEN_5606 : _GEN_5472; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5661 = _T_1007 ? _GEN_5607 : _GEN_5473; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5662 = _T_1007 ? _GEN_5608 : _GEN_5474; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5663 = _T_1007 ? _GEN_5609 : _GEN_5475; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5664 = _T_1007 ? _GEN_5610 : _GEN_5476; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5665 = _T_1007 ? _GEN_5611 : _GEN_5477; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5666 = _T_1007 ? _GEN_5612 : _GEN_5478; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5667 = _T_1007 ? _GEN_5613 : _GEN_5479; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5668 = _T_1007 ? _GEN_5614 : _GEN_5480; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5669 = _T_1007 ? _GEN_5615 : _GEN_5481; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5670 = _T_1007 ? _GEN_5616 : _GEN_5482; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5671 = _T_1007 ? _GEN_5617 : _GEN_5483; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5672 = _T_1007 ? _GEN_5618 : _GEN_5484; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5673 = _T_1007 ? _GEN_5619 : _GEN_5485; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5674 = _T_1007 ? _GEN_5620 : _GEN_5486; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5675 = _T_1007 ? _GEN_5621 : _GEN_5487; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5676 = _T_1007 ? _GEN_5622 : _GEN_5488; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5678 = _T_1007 ? _GEN_5624 : _GEN_5490; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [31:0] _GEN_5679 = _T_1007 ? _GEN_5625 : _GEN_5491; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [2:0] _funct3_T_71 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_1045 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _next_reg_has_T_108 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_109 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_110 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_111 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_112 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_113 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_114 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_115 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_116 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_117 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_118 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_119 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_120 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_121 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_122 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_123 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_124 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_125 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_126 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_127 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_128 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_129 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_130 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_131 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_132 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_133 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_134 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  next_reg_has_4 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_nowCSR_T_108 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_109 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_110 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_111 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_112 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_113 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_114 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_115 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_116 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_117 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_118 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_119 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_120 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_121 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_122 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_123 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_124 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_125 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_126 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_127 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_128 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_129 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_130 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_131 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_132 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_133 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_134 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] next_reg_nowCSR_4 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rmask_T_164 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_165 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_166 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_167 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_168 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_169 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_170 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_171 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_172 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_173 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_174 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_175 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_176 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_177 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _next_reg_rmask_T_178 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_179 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_180 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_181 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_182 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_183 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_184 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_185 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_186 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_187 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_188 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_189 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_190 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_191 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_192 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_193 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_194 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_195 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_196 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_197 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_198 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_199 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_200 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_201 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_202 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_203 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_204 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] next_reg_rmask_4 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_T_201 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] _next_reg_rData_T_24 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rData_T_25 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5682 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire  _next_reg_T_202 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_203 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _next_reg_rData_T_26 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _next_reg_rData_T_27 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _next_reg_rData_T_28 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _next_reg_rData_T_29 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [31:0] _GEN_5683 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5684 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_204 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] next_reg_rData_4 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5685 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_T_205 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_rd_46 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5686 = 5'h0 == rd ? rData_3 : _GEN_5638; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5687 = 5'h1 == rd ? rData_3 : _GEN_5639; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5688 = 5'h2 == rd ? rData_3 : _GEN_5640; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5689 = 5'h3 == rd ? rData_3 : _GEN_5641; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5690 = 5'h4 == rd ? rData_3 : _GEN_5642; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5691 = 5'h5 == rd ? rData_3 : _GEN_5643; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5692 = 5'h6 == rd ? rData_3 : _GEN_5644; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5693 = 5'h7 == rd ? rData_3 : _GEN_5645; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5694 = 5'h8 == rd ? rData_3 : _GEN_5646; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5695 = 5'h9 == rd ? rData_3 : _GEN_5647; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5696 = 5'ha == rd ? rData_3 : _GEN_5648; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5697 = 5'hb == rd ? rData_3 : _GEN_5649; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5698 = 5'hc == rd ? rData_3 : _GEN_5650; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5699 = 5'hd == rd ? rData_3 : _GEN_5651; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5700 = 5'he == rd ? rData_3 : _GEN_5652; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5701 = 5'hf == rd ? rData_3 : _GEN_5653; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5702 = 5'h10 == rd ? rData_3 : _GEN_5654; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5703 = 5'h11 == rd ? rData_3 : _GEN_5655; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5704 = 5'h12 == rd ? rData_3 : _GEN_5656; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5705 = 5'h13 == rd ? rData_3 : _GEN_5657; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5706 = 5'h14 == rd ? rData_3 : _GEN_5658; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5707 = 5'h15 == rd ? rData_3 : _GEN_5659; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5708 = 5'h16 == rd ? rData_3 : _GEN_5660; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5709 = 5'h17 == rd ? rData_3 : _GEN_5661; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5710 = 5'h18 == rd ? rData_3 : _GEN_5662; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5711 = 5'h19 == rd ? rData_3 : _GEN_5663; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5712 = 5'h1a == rd ? rData_3 : _GEN_5664; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5713 = 5'h1b == rd ? rData_3 : _GEN_5665; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5714 = 5'h1c == rd ? rData_3 : _GEN_5666; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5715 = 5'h1d == rd ? rData_3 : _GEN_5667; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5716 = 5'h1e == rd ? rData_3 : _GEN_5668; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [31:0] _GEN_5717 = 5'h1f == rd ? rData_3 : _GEN_5669; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire  _T_1054 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_1058 = csrAddr == 12'h301; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1059 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_misa_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_misa_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_misa_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5722 = csrAddr == 12'h301 ? _T_1057 : _GEN_5670; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1060 = csrAddr == 12'hf11; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1061 = csrAddr == 12'hf12; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1062 = csrAddr == 12'hf13; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1063 = csrAddr == 12'hf14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1064 = csrAddr == 12'h300; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1065 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_26 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_27 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mstatus_T_28 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mstatus_T_29 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_30 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mstatus_T_31 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mstatus_mstatusOld_WIRE_9 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire  next_csr_mstatus_mstatusOld_4_pad4 = _T_1057[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sie = _T_1057[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_pad3 = _T_1057[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mie = _T_1057[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_pad2 = _T_1057[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_spie = _T_1057[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_ube = _T_1057[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mpie = _T_1057[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_spp = _T_1057[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_vs = _T_1057[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_mpp = _T_1057[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_fs = _T_1057[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_xs = _T_1057[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mprv = _T_1057[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sum = _T_1057[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mxr = _T_1057[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_tvm = _T_1057[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_tw = _T_1057[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_tsr = _T_1057[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] next_csr_mstatus_mstatusOld_4_pad0 = _T_1057[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sd = _T_1057[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_8_fs = next_csr_mstatus_mstatusOld_4_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_95 = next_csr_mstatus_mstatusOld_4_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusNew_T_12 = next_csr_mstatus_mstatusOld_4_fs == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:42]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_sie = next_csr_mstatus_mstatusOld_4_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_85 = next_csr_mstatus_mstatusOld_4_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_pad4 = next_csr_mstatus_mstatusOld_4_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_84 = next_csr_mstatus_mstatusOld_4_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_lo_4 = {next_csr_mstatus_mstatusOld_4_sie,
    next_csr_mstatus_mstatusOld_4_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_pad2 = next_csr_mstatus_mstatusOld_4_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_88 = next_csr_mstatus_mstatusOld_4_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_mie = next_csr_mstatus_mstatusOld_4_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_87 = next_csr_mstatus_mstatusOld_4_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_pad2,
    next_csr_mstatus_mstatusOld_4_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_pad3 = next_csr_mstatus_mstatusOld_4_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_86 = next_csr_mstatus_mstatusOld_4_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_lo_hi_4 = {next_csr_mstatus_mstatusOld_4_pad2,
    next_csr_mstatus_mstatusOld_4_mie,next_csr_mstatus_mstatusOld_4_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [4:0] next_csr_mstatus_mstatusNew_lo_lo_4 = {next_csr_mstatus_mstatusOld_4_pad2,next_csr_mstatus_mstatusOld_4_mie
    ,next_csr_mstatus_mstatusOld_4_pad3,next_csr_mstatus_mstatusOld_4_sie,next_csr_mstatus_mstatusOld_4_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_ube = next_csr_mstatus_mstatusOld_4_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_90 = next_csr_mstatus_mstatusOld_4_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_spie = next_csr_mstatus_mstatusOld_4_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_89 = next_csr_mstatus_mstatusOld_4_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_hi_lo_4 = {next_csr_mstatus_mstatusOld_4_ube,
    next_csr_mstatus_mstatusOld_4_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_8_vs = next_csr_mstatus_mstatusOld_4_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_93 = next_csr_mstatus_mstatusOld_4_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_spp = next_csr_mstatus_mstatusOld_4_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_92 = next_csr_mstatus_mstatusOld_4_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_hi_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_vs,
    next_csr_mstatus_mstatusOld_4_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_mpie = next_csr_mstatus_mstatusOld_4_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_91 = next_csr_mstatus_mstatusOld_4_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_lo_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_vs,
    next_csr_mstatus_mstatusOld_4_spp,next_csr_mstatus_mstatusOld_4_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_hi_4 = {next_csr_mstatus_mstatusOld_4_vs,next_csr_mstatus_mstatusOld_4_spp,
    next_csr_mstatus_mstatusOld_4_mpie,next_csr_mstatus_mstatusOld_4_ube,next_csr_mstatus_mstatusOld_4_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [10:0] next_csr_mstatus_mstatusNew_lo_4 = {next_csr_mstatus_mstatusOld_4_vs,next_csr_mstatus_mstatusOld_4_spp,
    next_csr_mstatus_mstatusOld_4_mpie,next_csr_mstatus_mstatusOld_4_ube,next_csr_mstatus_mstatusOld_4_spie,
    next_csr_mstatus_mstatusOld_4_pad2,next_csr_mstatus_mstatusOld_4_mie,next_csr_mstatus_mstatusOld_4_pad3,
    next_csr_mstatus_mstatusOld_4_sie,next_csr_mstatus_mstatusOld_4_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_8_mpp = next_csr_mstatus_mstatusOld_4_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_94 = next_csr_mstatus_mstatusOld_4_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_lo_4 = {next_csr_mstatus_mstatusOld_4_fs,
    next_csr_mstatus_mstatusOld_4_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_sum = next_csr_mstatus_mstatusOld_4_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_98 = next_csr_mstatus_mstatusOld_4_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_mprv = next_csr_mstatus_mstatusOld_4_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_97 = next_csr_mstatus_mstatusOld_4_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_lo_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_sum,
    next_csr_mstatus_mstatusOld_4_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_8_xs = next_csr_mstatus_mstatusOld_4_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_96 = next_csr_mstatus_mstatusOld_4_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_hi_4 = {next_csr_mstatus_mstatusOld_4_sum,
    next_csr_mstatus_mstatusOld_4_mprv,next_csr_mstatus_mstatusOld_4_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [7:0] next_csr_mstatus_mstatusNew_hi_lo_4 = {next_csr_mstatus_mstatusOld_4_sum,next_csr_mstatus_mstatusOld_4_mprv
    ,next_csr_mstatus_mstatusOld_4_xs,next_csr_mstatus_mstatusOld_4_fs,next_csr_mstatus_mstatusOld_4_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_tw = next_csr_mstatus_mstatusOld_4_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_101 = next_csr_mstatus_mstatusOld_4_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_tvm = next_csr_mstatus_mstatusOld_4_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_100 = next_csr_mstatus_mstatusOld_4_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_hi_lo_hi_4 = {next_csr_mstatus_mstatusOld_4_tw,
    next_csr_mstatus_mstatusOld_4_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_mxr = next_csr_mstatus_mstatusOld_4_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_99 = next_csr_mstatus_mstatusOld_4_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_hi_hi_lo_4 = {next_csr_mstatus_mstatusOld_4_tw,
    next_csr_mstatus_mstatusOld_4_tvm,next_csr_mstatus_mstatusOld_4_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_sd = next_csr_mstatus_mstatusOld_4_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_104 = next_csr_mstatus_mstatusOld_4_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_WIRE_8_pad0 = next_csr_mstatus_mstatusOld_4_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_T_103 = next_csr_mstatus_mstatusOld_4_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusNew_hi_hi_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_sd,
    next_csr_mstatus_mstatusOld_4_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_8_tsr = next_csr_mstatus_mstatusOld_4_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_102 = next_csr_mstatus_mstatusOld_4_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [9:0] next_csr_mstatus_mstatusNew_hi_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_sd,
    next_csr_mstatus_mstatusOld_4_pad0,next_csr_mstatus_mstatusOld_4_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [12:0] next_csr_mstatus_mstatusNew_hi_hi_4 = {next_csr_mstatus_mstatusOld_4_sd,next_csr_mstatus_mstatusOld_4_pad0
    ,next_csr_mstatus_mstatusOld_4_tsr,next_csr_mstatus_mstatusOld_4_tw,next_csr_mstatus_mstatusOld_4_tvm,
    next_csr_mstatus_mstatusOld_4_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [20:0] next_csr_mstatus_mstatusNew_hi_4 = {next_csr_mstatus_mstatusOld_4_sd,next_csr_mstatus_mstatusOld_4_pad0,
    next_csr_mstatus_mstatusOld_4_tsr,next_csr_mstatus_mstatusOld_4_tw,next_csr_mstatus_mstatusOld_4_tvm,
    next_csr_mstatus_mstatusOld_4_mxr,next_csr_mstatus_mstatusNew_hi_lo_4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [31:0] _next_csr_mstatus_mstatusNew_T_13 = {next_csr_mstatus_mstatusOld_4_sd,next_csr_mstatus_mstatusOld_4_pad0,
    next_csr_mstatus_mstatusOld_4_tsr,next_csr_mstatus_mstatusOld_4_tw,next_csr_mstatus_mstatusOld_4_tvm,
    next_csr_mstatus_mstatusOld_4_mxr,next_csr_mstatus_mstatusNew_hi_lo_4,next_csr_mstatus_mstatusNew_lo_4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [30:0] _next_csr_mstatus_mstatusNew_T_14 = _next_csr_mstatus_mstatusNew_T_13[30:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:72]
  wire [31:0] next_csr_mstatus_mstatusNew_4 = {next_csr_mstatus_mstatusOld_4_fs == 2'h3,
    _next_csr_mstatus_mstatusNew_T_13[30:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [31:0] _GEN_5723 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_4 : _GEN_5671; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1066 = csrAddr == 12'h340; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1067 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mscratch_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mscratch_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mscratch_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5724 = csrAddr == 12'h340 ? _T_1057 : _GEN_5672; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1068 = csrAddr == 12'h305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1069 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtvec_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtvec_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mtvec_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5725 = csrAddr == 12'h305 ? _T_1057 : _GEN_5673; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1070 = csrAddr == 12'h306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1071 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcounteren_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcounteren_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mcounteren_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5726 = csrAddr == 12'h306 ? _T_1057 : _GEN_5674; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1072 = csrAddr == 12'h344; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [10:0] _next_csr_mip_T_16 = 11'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mip_T_17 = io_now_csr_mip & 32'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mip_T_18 = _T_1057 & 32'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [31:0] _next_csr_mip_T_19 = _next_csr_mip_T_1 | _next_csr_mip_T_18; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [31:0] _GEN_5727 = csrAddr == 12'h344 ? _next_csr_mip_T_19 : _GEN_5675; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1073 = csrAddr == 12'h304; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1074 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mie_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mie_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mie_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5728 = csrAddr == 12'h304 ? _T_1057 : _GEN_5676; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _T_1076 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire  _T_1077 = csrAddr == 12'h342; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1078 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_24 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_25 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcause_T_26 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcause_T_27 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_28 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mcause_T_29 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5730 = csrAddr == 12'h342 ? _T_1057 : _GEN_5678; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1079 = csrAddr == 12'h343; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1080 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_42 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_43 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtval_T_44 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtval_T_45 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_46 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _next_csr_mtval_T_47 = rData_3 | _T_1096; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [31:0] _GEN_5731 = csrAddr == 12'h343 ? _T_1057 : _GEN_5679; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5732 = has_15 ? _GEN_5722 : _GEN_5670; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5733 = has_15 ? _GEN_5723 : _GEN_5671; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5734 = has_15 ? _GEN_5724 : _GEN_5672; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5735 = has_15 ? _GEN_5725 : _GEN_5673; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5736 = has_15 ? _GEN_5726 : _GEN_5674; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5737 = has_15 ? _GEN_5727 : _GEN_5675; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5738 = has_15 ? _GEN_5728 : _GEN_5676; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5740 = has_15 ? _GEN_5730 : _GEN_5678; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5741 = has_15 ? _GEN_5731 : _GEN_5679; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5744 = _T_1090 ? _GEN_5732 : _GEN_5670; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5745 = _T_1090 ? _GEN_5733 : _GEN_5671; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5746 = _T_1090 ? _GEN_5734 : _GEN_5672; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5747 = _T_1090 ? _GEN_5735 : _GEN_5673; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5748 = _T_1090 ? _GEN_5736 : _GEN_5674; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5749 = _T_1090 ? _GEN_5737 : _GEN_5675; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5750 = _T_1090 ? _GEN_5738 : _GEN_5676; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5752 = _T_1090 ? _GEN_5740 : _GEN_5678; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5753 = _T_1090 ? _GEN_5741 : _GEN_5679; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [31:0] _GEN_5756 = ~isIllegalWrite_4 ? _GEN_5686 : _GEN_5638; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5757 = ~isIllegalWrite_4 ? _GEN_5687 : _GEN_5639; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5758 = ~isIllegalWrite_4 ? _GEN_5688 : _GEN_5640; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5759 = ~isIllegalWrite_4 ? _GEN_5689 : _GEN_5641; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5760 = ~isIllegalWrite_4 ? _GEN_5690 : _GEN_5642; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5761 = ~isIllegalWrite_4 ? _GEN_5691 : _GEN_5643; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5762 = ~isIllegalWrite_4 ? _GEN_5692 : _GEN_5644; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5763 = ~isIllegalWrite_4 ? _GEN_5693 : _GEN_5645; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5764 = ~isIllegalWrite_4 ? _GEN_5694 : _GEN_5646; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5765 = ~isIllegalWrite_4 ? _GEN_5695 : _GEN_5647; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5766 = ~isIllegalWrite_4 ? _GEN_5696 : _GEN_5648; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5767 = ~isIllegalWrite_4 ? _GEN_5697 : _GEN_5649; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5768 = ~isIllegalWrite_4 ? _GEN_5698 : _GEN_5650; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5769 = ~isIllegalWrite_4 ? _GEN_5699 : _GEN_5651; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5770 = ~isIllegalWrite_4 ? _GEN_5700 : _GEN_5652; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5771 = ~isIllegalWrite_4 ? _GEN_5701 : _GEN_5653; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5772 = ~isIllegalWrite_4 ? _GEN_5702 : _GEN_5654; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5773 = ~isIllegalWrite_4 ? _GEN_5703 : _GEN_5655; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5774 = ~isIllegalWrite_4 ? _GEN_5704 : _GEN_5656; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5775 = ~isIllegalWrite_4 ? _GEN_5705 : _GEN_5657; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5776 = ~isIllegalWrite_4 ? _GEN_5706 : _GEN_5658; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5777 = ~isIllegalWrite_4 ? _GEN_5707 : _GEN_5659; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5778 = ~isIllegalWrite_4 ? _GEN_5708 : _GEN_5660; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5779 = ~isIllegalWrite_4 ? _GEN_5709 : _GEN_5661; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5780 = ~isIllegalWrite_4 ? _GEN_5710 : _GEN_5662; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5781 = ~isIllegalWrite_4 ? _GEN_5711 : _GEN_5663; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5782 = ~isIllegalWrite_4 ? _GEN_5712 : _GEN_5664; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5783 = ~isIllegalWrite_4 ? _GEN_5713 : _GEN_5665; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5784 = ~isIllegalWrite_4 ? _GEN_5714 : _GEN_5666; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5785 = ~isIllegalWrite_4 ? _GEN_5715 : _GEN_5667; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5786 = ~isIllegalWrite_4 ? _GEN_5716 : _GEN_5668; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5787 = ~isIllegalWrite_4 ? _GEN_5717 : _GEN_5669; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5788 = ~isIllegalWrite_4 ? _GEN_5744 : _GEN_5670; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5789 = ~isIllegalWrite_4 ? _GEN_5745 : _GEN_5671; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5790 = ~isIllegalWrite_4 ? _GEN_5746 : _GEN_5672; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5791 = ~isIllegalWrite_4 ? _GEN_5747 : _GEN_5673; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5792 = ~isIllegalWrite_4 ? _GEN_5748 : _GEN_5674; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5793 = ~isIllegalWrite_4 ? _GEN_5749 : _GEN_5675; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5794 = ~isIllegalWrite_4 ? _GEN_5750 : _GEN_5676; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5796 = ~isIllegalWrite_4 ? _GEN_5752 : _GEN_5678; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [31:0] _GEN_5797 = ~isIllegalWrite_4 ? _GEN_5753 : _GEN_5679; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [2:0] _GEN_5803 = _T_1041 ? inst[14:12] : _GEN_5631; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5805 = _T_1041 ? inst[6:0] : _GEN_5633; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_5810 = _T_1041 ? _GEN_5756 : _GEN_5638; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5811 = _T_1041 ? _GEN_5757 : _GEN_5639; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5812 = _T_1041 ? _GEN_5758 : _GEN_5640; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5813 = _T_1041 ? _GEN_5759 : _GEN_5641; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5814 = _T_1041 ? _GEN_5760 : _GEN_5642; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5815 = _T_1041 ? _GEN_5761 : _GEN_5643; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5816 = _T_1041 ? _GEN_5762 : _GEN_5644; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5817 = _T_1041 ? _GEN_5763 : _GEN_5645; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5818 = _T_1041 ? _GEN_5764 : _GEN_5646; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5819 = _T_1041 ? _GEN_5765 : _GEN_5647; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5820 = _T_1041 ? _GEN_5766 : _GEN_5648; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5821 = _T_1041 ? _GEN_5767 : _GEN_5649; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5822 = _T_1041 ? _GEN_5768 : _GEN_5650; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5823 = _T_1041 ? _GEN_5769 : _GEN_5651; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5824 = _T_1041 ? _GEN_5770 : _GEN_5652; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5825 = _T_1041 ? _GEN_5771 : _GEN_5653; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5826 = _T_1041 ? _GEN_5772 : _GEN_5654; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5827 = _T_1041 ? _GEN_5773 : _GEN_5655; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5828 = _T_1041 ? _GEN_5774 : _GEN_5656; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5829 = _T_1041 ? _GEN_5775 : _GEN_5657; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5830 = _T_1041 ? _GEN_5776 : _GEN_5658; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5831 = _T_1041 ? _GEN_5777 : _GEN_5659; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5832 = _T_1041 ? _GEN_5778 : _GEN_5660; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5833 = _T_1041 ? _GEN_5779 : _GEN_5661; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5834 = _T_1041 ? _GEN_5780 : _GEN_5662; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5835 = _T_1041 ? _GEN_5781 : _GEN_5663; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5836 = _T_1041 ? _GEN_5782 : _GEN_5664; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5837 = _T_1041 ? _GEN_5783 : _GEN_5665; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5838 = _T_1041 ? _GEN_5784 : _GEN_5666; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5839 = _T_1041 ? _GEN_5785 : _GEN_5667; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5840 = _T_1041 ? _GEN_5786 : _GEN_5668; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5841 = _T_1041 ? _GEN_5787 : _GEN_5669; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5842 = _T_1041 ? _GEN_5788 : _GEN_5670; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5843 = _T_1041 ? _GEN_5789 : _GEN_5671; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5844 = _T_1041 ? _GEN_5790 : _GEN_5672; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5845 = _T_1041 ? _GEN_5791 : _GEN_5673; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5846 = _T_1041 ? _GEN_5792 : _GEN_5674; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5847 = _T_1041 ? _GEN_5793 : _GEN_5675; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5848 = _T_1041 ? _GEN_5794 : _GEN_5676; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5850 = _T_1041 ? _GEN_5796 : _GEN_5678; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [31:0] _GEN_5851 = _T_1041 ? _GEN_5797 : _GEN_5679; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [2:0] _funct3_T_72 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_1086 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _next_reg_has_T_135 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_136 = _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_137 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_138 = _has_T_407 | _has_T_405; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_139 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_140 = _has_T_409 | _has_T_408; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_141 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_142 = _has_T_411 | _has_T_410; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_143 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_144 = _has_T_413 | _has_T_412; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_145 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_146 = _has_T_415 | _has_T_414; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_147 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_148 = _has_T_417 | _has_T_416; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_149 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_150 = _has_T_419 | _has_T_418; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_151 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_152 = _has_T_421 | _has_T_420; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_153 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_154 = _has_T_423 | _has_T_422; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_155 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_156 = _has_T_425 | _has_T_424; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_157 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_158 = _has_T_427 | _has_T_426; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_159 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_160 = _has_T_429 | _has_T_428; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_has_T_161 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  next_reg_has_5 = _has_T_431 | _has_T_430; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 23:48]
  wire  _next_reg_nowCSR_T_135 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_136 = _has_T_405 ? io_now_csr_misa : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_137 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_138 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_139 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_140 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_141 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_142 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_143 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_144 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_145 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_146 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_147 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_148 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_149 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_150 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_151 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_152 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_153 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_154 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_155 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_156 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_157 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_158 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_159 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_nowCSR_T_160 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire  _next_reg_nowCSR_T_161 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] next_reg_nowCSR_5 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rmask_T_205 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_206 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_207 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_208 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_209 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_210 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_211 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_212 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_213 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_214 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_215 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_216 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_217 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire [31:0] _next_reg_rmask_T_218 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 29:40]
  wire  _next_reg_rmask_T_219 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_220 = _has_T_405 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_221 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_222 = _has_T_407 ? 32'hffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_223 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_224 = _has_T_409 ? 32'hffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_225 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_226 = _has_T_411 ? 32'hffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_227 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_228 = _has_T_413 ? 32'hffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_229 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_230 = _has_T_415 ? 32'hffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_231 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_232 = _has_T_417 ? 32'hffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_233 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_234 = _has_T_419 ? 32'hffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_235 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_236 = _has_T_421 ? 32'hffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_237 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_238 = _has_T_423 ? 32'hffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_239 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_240 = _has_T_425 ? 32'hffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_241 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_242 = _has_T_427 ? 32'hffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_243 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] _next_reg_rmask_T_244 = _has_T_429 ? 32'hffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_rmask_T_245 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [31:0] next_reg_rmask_5 = _has_T_431 ? 32'hffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire  _next_reg_T_206 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] _next_reg_rData_T_30 = nowCSR_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [31:0] _next_reg_rData_T_31 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [31:0] _GEN_5854 = has_15 ? _rData_T_19 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire  _next_reg_T_207 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_208 = io_now_csr_IALIGN == 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:31]
  wire [29:0] _next_reg_rData_T_32 = 30'h3fffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:30]
  wire [31:0] _next_reg_rData_T_33 = 32'hfffffffc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:25]
  wire [31:0] _next_reg_rData_T_34 = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:77]
  wire [31:0] _next_reg_rData_T_35 = 32'hfffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [31:0] _GEN_5855 = io_now_csr_IALIGN == 8'h20 ? _rData_T_23 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [31:0] _GEN_5856 = _has_T_427 ? _GEN_5891 : _GEN_5890; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire  _next_reg_T_209 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [31:0] next_reg_rData_5 = _T_1123 ? _GEN_5892 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5857 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_T_210 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _next_reg_rd_47 = rData_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [31:0] _GEN_5858 = 5'h0 == rd ? rData_3 : _GEN_5810; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5859 = 5'h1 == rd ? rData_3 : _GEN_5811; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5860 = 5'h2 == rd ? rData_3 : _GEN_5812; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5861 = 5'h3 == rd ? rData_3 : _GEN_5813; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5862 = 5'h4 == rd ? rData_3 : _GEN_5814; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5863 = 5'h5 == rd ? rData_3 : _GEN_5815; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5864 = 5'h6 == rd ? rData_3 : _GEN_5816; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5865 = 5'h7 == rd ? rData_3 : _GEN_5817; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5866 = 5'h8 == rd ? rData_3 : _GEN_5818; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5867 = 5'h9 == rd ? rData_3 : _GEN_5819; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5868 = 5'ha == rd ? rData_3 : _GEN_5820; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5869 = 5'hb == rd ? rData_3 : _GEN_5821; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5870 = 5'hc == rd ? rData_3 : _GEN_5822; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5871 = 5'hd == rd ? rData_3 : _GEN_5823; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5872 = 5'he == rd ? rData_3 : _GEN_5824; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5873 = 5'hf == rd ? rData_3 : _GEN_5825; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5874 = 5'h10 == rd ? rData_3 : _GEN_5826; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5875 = 5'h11 == rd ? rData_3 : _GEN_5827; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5876 = 5'h12 == rd ? rData_3 : _GEN_5828; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5877 = 5'h13 == rd ? rData_3 : _GEN_5829; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5878 = 5'h14 == rd ? rData_3 : _GEN_5830; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5879 = 5'h15 == rd ? rData_3 : _GEN_5831; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5880 = 5'h16 == rd ? rData_3 : _GEN_5832; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5881 = 5'h17 == rd ? rData_3 : _GEN_5833; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5882 = 5'h18 == rd ? rData_3 : _GEN_5834; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5883 = 5'h19 == rd ? rData_3 : _GEN_5835; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5884 = 5'h1a == rd ? rData_3 : _GEN_5836; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5885 = 5'h1b == rd ? rData_3 : _GEN_5837; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5886 = 5'h1c == rd ? rData_3 : _GEN_5838; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5887 = 5'h1d == rd ? rData_3 : _GEN_5839; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5888 = 5'h1e == rd ? rData_3 : _GEN_5840; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [31:0] _GEN_5889 = 5'h1f == rd ? rData_3 : _GEN_5841; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire  _T_1094 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire  _T_1099 = csrAddr == 12'h301; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1100 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_misa_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_misa_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_misa_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_misa_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5894 = csrAddr == 12'h301 ? _T_1098 : _GEN_5842; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1101 = csrAddr == 12'hf11; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1102 = csrAddr == 12'hf12; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1103 = csrAddr == 12'hf13; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1104 = csrAddr == 12'hf14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire  _T_1105 = csrAddr == 12'h300; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1106 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_32 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_33 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mstatus_T_34 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mstatus_T_35 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mstatus_T_36 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mstatus_T_37 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mstatus_mstatusOld_WIRE_11 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire  next_csr_mstatus_mstatusOld_5_pad4 = _T_1098[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sie = _T_1098[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_pad3 = _T_1098[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mie = _T_1098[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_pad2 = _T_1098[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_spie = _T_1098[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_ube = _T_1098[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mpie = _T_1098[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_spp = _T_1098[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_vs = _T_1098[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_mpp = _T_1098[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_fs = _T_1098[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_xs = _T_1098[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mprv = _T_1098[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sum = _T_1098[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mxr = _T_1098[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_tvm = _T_1098[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_tw = _T_1098[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_tsr = _T_1098[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] next_csr_mstatus_mstatusOld_5_pad0 = _T_1098[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sd = _T_1098[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_10_fs = next_csr_mstatus_mstatusOld_5_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_116 = next_csr_mstatus_mstatusOld_5_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusNew_T_15 = next_csr_mstatus_mstatusOld_5_fs == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:42]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_sie = next_csr_mstatus_mstatusOld_5_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_106 = next_csr_mstatus_mstatusOld_5_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_pad4 = next_csr_mstatus_mstatusOld_5_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_105 = next_csr_mstatus_mstatusOld_5_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_lo_5 = {next_csr_mstatus_mstatusOld_5_sie,
    next_csr_mstatus_mstatusOld_5_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_pad2 = next_csr_mstatus_mstatusOld_5_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_109 = next_csr_mstatus_mstatusOld_5_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_mie = next_csr_mstatus_mstatusOld_5_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_108 = next_csr_mstatus_mstatusOld_5_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_lo_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_pad2,
    next_csr_mstatus_mstatusOld_5_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_pad3 = next_csr_mstatus_mstatusOld_5_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_107 = next_csr_mstatus_mstatusOld_5_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_lo_hi_5 = {next_csr_mstatus_mstatusOld_5_pad2,
    next_csr_mstatus_mstatusOld_5_mie,next_csr_mstatus_mstatusOld_5_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [4:0] next_csr_mstatus_mstatusNew_lo_lo_5 = {next_csr_mstatus_mstatusOld_5_pad2,next_csr_mstatus_mstatusOld_5_mie
    ,next_csr_mstatus_mstatusOld_5_pad3,next_csr_mstatus_mstatusOld_5_sie,next_csr_mstatus_mstatusOld_5_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_ube = next_csr_mstatus_mstatusOld_5_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_111 = next_csr_mstatus_mstatusOld_5_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_spie = next_csr_mstatus_mstatusOld_5_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_110 = next_csr_mstatus_mstatusOld_5_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_lo_hi_lo_5 = {next_csr_mstatus_mstatusOld_5_ube,
    next_csr_mstatus_mstatusOld_5_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_10_vs = next_csr_mstatus_mstatusOld_5_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_114 = next_csr_mstatus_mstatusOld_5_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_spp = next_csr_mstatus_mstatusOld_5_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_113 = next_csr_mstatus_mstatusOld_5_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_lo_hi_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_vs,
    next_csr_mstatus_mstatusOld_5_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_mpie = next_csr_mstatus_mstatusOld_5_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_112 = next_csr_mstatus_mstatusOld_5_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_lo_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_vs,
    next_csr_mstatus_mstatusOld_5_spp,next_csr_mstatus_mstatusOld_5_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_hi_5 = {next_csr_mstatus_mstatusOld_5_vs,next_csr_mstatus_mstatusOld_5_spp,
    next_csr_mstatus_mstatusOld_5_mpie,next_csr_mstatus_mstatusOld_5_ube,next_csr_mstatus_mstatusOld_5_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [10:0] next_csr_mstatus_mstatusNew_lo_5 = {next_csr_mstatus_mstatusOld_5_vs,next_csr_mstatus_mstatusOld_5_spp,
    next_csr_mstatus_mstatusOld_5_mpie,next_csr_mstatus_mstatusOld_5_ube,next_csr_mstatus_mstatusOld_5_spie,
    next_csr_mstatus_mstatusOld_5_pad2,next_csr_mstatus_mstatusOld_5_mie,next_csr_mstatus_mstatusOld_5_pad3,
    next_csr_mstatus_mstatusOld_5_sie,next_csr_mstatus_mstatusOld_5_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_10_mpp = next_csr_mstatus_mstatusOld_5_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_115 = next_csr_mstatus_mstatusOld_5_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_lo_5 = {next_csr_mstatus_mstatusOld_5_fs,
    next_csr_mstatus_mstatusOld_5_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_sum = next_csr_mstatus_mstatusOld_5_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_119 = next_csr_mstatus_mstatusOld_5_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_mprv = next_csr_mstatus_mstatusOld_5_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_118 = next_csr_mstatus_mstatusOld_5_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_lo_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_sum,
    next_csr_mstatus_mstatusOld_5_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [1:0] _next_csr_mstatus_mstatusOld_WIRE_10_xs = next_csr_mstatus_mstatusOld_5_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] _next_csr_mstatus_mstatusOld_T_117 = next_csr_mstatus_mstatusOld_5_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [3:0] next_csr_mstatus_mstatusNew_hi_lo_hi_5 = {next_csr_mstatus_mstatusOld_5_sum,
    next_csr_mstatus_mstatusOld_5_mprv,next_csr_mstatus_mstatusOld_5_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [7:0] next_csr_mstatus_mstatusNew_hi_lo_5 = {next_csr_mstatus_mstatusOld_5_sum,next_csr_mstatus_mstatusOld_5_mprv
    ,next_csr_mstatus_mstatusOld_5_xs,next_csr_mstatus_mstatusOld_5_fs,next_csr_mstatus_mstatusOld_5_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_tw = next_csr_mstatus_mstatusOld_5_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_122 = next_csr_mstatus_mstatusOld_5_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_tvm = next_csr_mstatus_mstatusOld_5_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_121 = next_csr_mstatus_mstatusOld_5_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusNew_hi_hi_lo_hi_5 = {next_csr_mstatus_mstatusOld_5_tw,
    next_csr_mstatus_mstatusOld_5_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_mxr = next_csr_mstatus_mstatusOld_5_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_120 = next_csr_mstatus_mstatusOld_5_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [2:0] next_csr_mstatus_mstatusNew_hi_hi_lo_5 = {next_csr_mstatus_mstatusOld_5_tw,
    next_csr_mstatus_mstatusOld_5_tvm,next_csr_mstatus_mstatusOld_5_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_sd = next_csr_mstatus_mstatusOld_5_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_125 = next_csr_mstatus_mstatusOld_5_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_WIRE_10_pad0 = next_csr_mstatus_mstatusOld_5_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [7:0] _next_csr_mstatus_mstatusOld_T_124 = next_csr_mstatus_mstatusOld_5_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusNew_hi_hi_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_sd,
    next_csr_mstatus_mstatusOld_5_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire  _next_csr_mstatus_mstatusOld_WIRE_10_tsr = next_csr_mstatus_mstatusOld_5_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  _next_csr_mstatus_mstatusOld_T_123 = next_csr_mstatus_mstatusOld_5_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [9:0] next_csr_mstatus_mstatusNew_hi_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_sd,
    next_csr_mstatus_mstatusOld_5_pad0,next_csr_mstatus_mstatusOld_5_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [12:0] next_csr_mstatus_mstatusNew_hi_hi_5 = {next_csr_mstatus_mstatusOld_5_sd,next_csr_mstatus_mstatusOld_5_pad0
    ,next_csr_mstatus_mstatusOld_5_tsr,next_csr_mstatus_mstatusOld_5_tw,next_csr_mstatus_mstatusOld_5_tvm,
    next_csr_mstatus_mstatusOld_5_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [20:0] next_csr_mstatus_mstatusNew_hi_5 = {next_csr_mstatus_mstatusOld_5_sd,next_csr_mstatus_mstatusOld_5_pad0,
    next_csr_mstatus_mstatusOld_5_tsr,next_csr_mstatus_mstatusOld_5_tw,next_csr_mstatus_mstatusOld_5_tvm,
    next_csr_mstatus_mstatusOld_5_mxr,next_csr_mstatus_mstatusNew_hi_lo_5}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [31:0] _next_csr_mstatus_mstatusNew_T_16 = {next_csr_mstatus_mstatusOld_5_sd,next_csr_mstatus_mstatusOld_5_pad0,
    next_csr_mstatus_mstatusOld_5_tsr,next_csr_mstatus_mstatusOld_5_tw,next_csr_mstatus_mstatusOld_5_tvm,
    next_csr_mstatus_mstatusOld_5_mxr,next_csr_mstatus_mstatusNew_hi_lo_5,next_csr_mstatus_mstatusNew_lo_5}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [30:0] _next_csr_mstatus_mstatusNew_T_17 = _next_csr_mstatus_mstatusNew_T_16[30:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:72]
  wire [31:0] next_csr_mstatus_mstatusNew_5 = {next_csr_mstatus_mstatusOld_5_fs == 2'h3,
    _next_csr_mstatus_mstatusNew_T_16[30:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [31:0] _GEN_5895 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_5 : _GEN_5843; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1107 = csrAddr == 12'h340; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1108 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mscratch_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mscratch_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mscratch_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mscratch_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5896 = csrAddr == 12'h340 ? _T_1098 : _GEN_5844; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1109 = csrAddr == 12'h305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1110 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtvec_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtvec_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtvec_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mtvec_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5897 = csrAddr == 12'h305 ? _T_1098 : _GEN_5845; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1111 = csrAddr == 12'h306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1112 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcounteren_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcounteren_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcounteren_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mcounteren_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5898 = csrAddr == 12'h306 ? _T_1098 : _GEN_5846; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1113 = csrAddr == 12'h344; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [10:0] _next_csr_mip_T_20 = 11'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mip_T_21 = io_now_csr_mip & 32'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mip_T_22 = _T_1098 & 32'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [31:0] _next_csr_mip_T_23 = _next_csr_mip_T_1 | _next_csr_mip_T_22; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [31:0] _GEN_5899 = csrAddr == 12'h344 ? _next_csr_mip_T_23 : _GEN_5847; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1114 = csrAddr == 12'h304; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1115 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mie_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mie_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mie_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mie_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5900 = csrAddr == 12'h304 ? _T_1098 : _GEN_5848; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _T_1117 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire  _T_1118 = csrAddr == 12'h342; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1119 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_30 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_31 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mcause_T_32 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mcause_T_33 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mcause_T_34 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mcause_T_35 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5902 = csrAddr == 12'h342 ? _T_1098 : _GEN_5850; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  _T_1120 = csrAddr == 12'h343; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:19]
  wire [31:0] _T_1121 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_48 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_49 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:53]
  wire [31:0] _next_csr_mtval_T_50 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [31:0] _next_csr_mtval_T_51 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 30:40]
  wire [31:0] _next_csr_mtval_T_52 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _next_csr_mtval_T_53 = rData_3 & _T_1097; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [31:0] _GEN_5903 = csrAddr == 12'h343 ? _T_1098 : _GEN_5851; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [31:0] _GEN_5904 = has_15 ? _GEN_5894 : _GEN_5842; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5905 = has_15 ? _GEN_5895 : _GEN_5843; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5906 = has_15 ? _GEN_5896 : _GEN_5844; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5907 = has_15 ? _GEN_5897 : _GEN_5845; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5908 = has_15 ? _GEN_5898 : _GEN_5846; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5909 = has_15 ? _GEN_5899 : _GEN_5847; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5910 = has_15 ? _GEN_5900 : _GEN_5848; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5912 = has_15 ? _GEN_5902 : _GEN_5850; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5913 = has_15 ? _GEN_5903 : _GEN_5851; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [31:0] _GEN_5916 = rs1 != 5'h0 ? _GEN_5904 : _GEN_5842; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5917 = rs1 != 5'h0 ? _GEN_5905 : _GEN_5843; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5918 = rs1 != 5'h0 ? _GEN_5906 : _GEN_5844; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5919 = rs1 != 5'h0 ? _GEN_5907 : _GEN_5845; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5920 = rs1 != 5'h0 ? _GEN_5908 : _GEN_5846; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5921 = rs1 != 5'h0 ? _GEN_5909 : _GEN_5847; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5922 = rs1 != 5'h0 ? _GEN_5910 : _GEN_5848; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5924 = rs1 != 5'h0 ? _GEN_5912 : _GEN_5850; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5925 = rs1 != 5'h0 ? _GEN_5913 : _GEN_5851; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [31:0] _GEN_5928 = ~isIllegalWrite_5 ? _GEN_5858 : _GEN_5810; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5929 = ~isIllegalWrite_5 ? _GEN_5859 : _GEN_5811; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5930 = ~isIllegalWrite_5 ? _GEN_5860 : _GEN_5812; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5931 = ~isIllegalWrite_5 ? _GEN_5861 : _GEN_5813; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5932 = ~isIllegalWrite_5 ? _GEN_5862 : _GEN_5814; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5933 = ~isIllegalWrite_5 ? _GEN_5863 : _GEN_5815; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5934 = ~isIllegalWrite_5 ? _GEN_5864 : _GEN_5816; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5935 = ~isIllegalWrite_5 ? _GEN_5865 : _GEN_5817; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5936 = ~isIllegalWrite_5 ? _GEN_5866 : _GEN_5818; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5937 = ~isIllegalWrite_5 ? _GEN_5867 : _GEN_5819; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5938 = ~isIllegalWrite_5 ? _GEN_5868 : _GEN_5820; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5939 = ~isIllegalWrite_5 ? _GEN_5869 : _GEN_5821; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5940 = ~isIllegalWrite_5 ? _GEN_5870 : _GEN_5822; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5941 = ~isIllegalWrite_5 ? _GEN_5871 : _GEN_5823; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5942 = ~isIllegalWrite_5 ? _GEN_5872 : _GEN_5824; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5943 = ~isIllegalWrite_5 ? _GEN_5873 : _GEN_5825; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5944 = ~isIllegalWrite_5 ? _GEN_5874 : _GEN_5826; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5945 = ~isIllegalWrite_5 ? _GEN_5875 : _GEN_5827; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5946 = ~isIllegalWrite_5 ? _GEN_5876 : _GEN_5828; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5947 = ~isIllegalWrite_5 ? _GEN_5877 : _GEN_5829; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5948 = ~isIllegalWrite_5 ? _GEN_5878 : _GEN_5830; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5949 = ~isIllegalWrite_5 ? _GEN_5879 : _GEN_5831; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5950 = ~isIllegalWrite_5 ? _GEN_5880 : _GEN_5832; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5951 = ~isIllegalWrite_5 ? _GEN_5881 : _GEN_5833; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5952 = ~isIllegalWrite_5 ? _GEN_5882 : _GEN_5834; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5953 = ~isIllegalWrite_5 ? _GEN_5883 : _GEN_5835; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5954 = ~isIllegalWrite_5 ? _GEN_5884 : _GEN_5836; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5955 = ~isIllegalWrite_5 ? _GEN_5885 : _GEN_5837; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5956 = ~isIllegalWrite_5 ? _GEN_5886 : _GEN_5838; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5957 = ~isIllegalWrite_5 ? _GEN_5887 : _GEN_5839; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5958 = ~isIllegalWrite_5 ? _GEN_5888 : _GEN_5840; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5959 = ~isIllegalWrite_5 ? _GEN_5889 : _GEN_5841; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5960 = ~isIllegalWrite_5 ? _GEN_5916 : _GEN_5842; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5961 = ~isIllegalWrite_5 ? _GEN_5917 : _GEN_5843; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5962 = ~isIllegalWrite_5 ? _GEN_5918 : _GEN_5844; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5963 = ~isIllegalWrite_5 ? _GEN_5919 : _GEN_5845; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5964 = ~isIllegalWrite_5 ? _GEN_5920 : _GEN_5846; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5965 = ~isIllegalWrite_5 ? _GEN_5921 : _GEN_5847; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5966 = ~isIllegalWrite_5 ? _GEN_5922 : _GEN_5848; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5968 = ~isIllegalWrite_5 ? _GEN_5924 : _GEN_5850; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [31:0] _GEN_5969 = ~isIllegalWrite_5 ? _GEN_5925 : _GEN_5851; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [2:0] _GEN_5975 = _T_1082 ? inst[14:12] : _GEN_5803; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5977 = _T_1082 ? inst[6:0] : _GEN_5805; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_5982 = _T_1082 ? _GEN_5928 : _GEN_5810; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5983 = _T_1082 ? _GEN_5929 : _GEN_5811; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5984 = _T_1082 ? _GEN_5930 : _GEN_5812; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5985 = _T_1082 ? _GEN_5931 : _GEN_5813; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5986 = _T_1082 ? _GEN_5932 : _GEN_5814; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5987 = _T_1082 ? _GEN_5933 : _GEN_5815; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5988 = _T_1082 ? _GEN_5934 : _GEN_5816; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5989 = _T_1082 ? _GEN_5935 : _GEN_5817; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5990 = _T_1082 ? _GEN_5936 : _GEN_5818; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5991 = _T_1082 ? _GEN_5937 : _GEN_5819; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5992 = _T_1082 ? _GEN_5938 : _GEN_5820; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5993 = _T_1082 ? _GEN_5939 : _GEN_5821; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5994 = _T_1082 ? _GEN_5940 : _GEN_5822; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5995 = _T_1082 ? _GEN_5941 : _GEN_5823; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5996 = _T_1082 ? _GEN_5942 : _GEN_5824; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5997 = _T_1082 ? _GEN_5943 : _GEN_5825; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5998 = _T_1082 ? _GEN_5944 : _GEN_5826; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_5999 = _T_1082 ? _GEN_5945 : _GEN_5827; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6000 = _T_1082 ? _GEN_5946 : _GEN_5828; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6001 = _T_1082 ? _GEN_5947 : _GEN_5829; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6002 = _T_1082 ? _GEN_5948 : _GEN_5830; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6003 = _T_1082 ? _GEN_5949 : _GEN_5831; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6004 = _T_1082 ? _GEN_5950 : _GEN_5832; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6005 = _T_1082 ? _GEN_5951 : _GEN_5833; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6006 = _T_1082 ? _GEN_5952 : _GEN_5834; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6007 = _T_1082 ? _GEN_5953 : _GEN_5835; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6008 = _T_1082 ? _GEN_5954 : _GEN_5836; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6009 = _T_1082 ? _GEN_5955 : _GEN_5837; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6010 = _T_1082 ? _GEN_5956 : _GEN_5838; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6011 = _T_1082 ? _GEN_5957 : _GEN_5839; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6012 = _T_1082 ? _GEN_5958 : _GEN_5840; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6013 = _T_1082 ? _GEN_5959 : _GEN_5841; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6014 = _T_1082 ? _GEN_5960 : _GEN_5842; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6015 = _T_1082 ? _GEN_5961 : _GEN_5843; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6016 = _T_1082 ? _GEN_5962 : _GEN_5844; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6017 = _T_1082 ? _GEN_5963 : _GEN_5845; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6018 = _T_1082 ? _GEN_5964 : _GEN_5846; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6019 = _T_1082 ? _GEN_5965 : _GEN_5847; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6020 = _T_1082 ? _GEN_5966 : _GEN_5848; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6022 = _T_1082 ? _GEN_5968 : _GEN_5850; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] _GEN_6023 = _T_1082 ? _GEN_5969 : _GEN_5851; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [31:0] now_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [1:0] _T_1137 = io_now_csr_stvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:27]
  wire  _T_1138 = 2'h0 == io_now_csr_stvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35]
  wire  _T_1139 = 2'h1 == io_now_csr_stvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35]
  wire  _GEN_6036 = 2'h1 == io_now_csr_stvec[1:0] | _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 316:29]
  wire  _GEN_6038 = 2'h0 == io_now_csr_stvec[1:0] | _GEN_6036; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 311:29]
  wire  _GEN_6048 = 8'h20 == io_now_csr_MXLEN ? _GEN_6038 : _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [1:0] _T_1153 = io_now_csr_mtvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:27]
  wire  _T_1154 = 2'h0 == io_now_csr_mtvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35]
  wire  _T_1155 = 2'h1 == io_now_csr_mtvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35]
  wire  _GEN_6056 = 2'h1 == io_now_csr_mtvec[1:0] | _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 242:29]
  wire  _GEN_6058 = 2'h0 == io_now_csr_mtvec[1:0] | _GEN_6056; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 237:29]
  wire  _GEN_6068 = _T_1123 ? _GEN_6058 : _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire  _GEN_6079 = delegS ? _GEN_6048 : _GEN_6068; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire  _GEN_6096 = raiseExceptionIntr ? _GEN_6079 : _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire  global_data_setpc = io_valid & _GEN_6096; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 113:21]
  wire  _GEN_6150 = global_data_setpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 113:21]
  wire  _T_1122 = ~global_data_setpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 150:10]
  wire [1:0] _next_pc_T_30 = inst[1:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:37]
  wire  _next_pc_T_31 = inst[1:0] == 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:44]
  wire [2:0] _next_pc_T_32 = inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:32]
  wire [31:0] _GEN_6214 = {{29'd0}, _next_pc_T_32}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [32:0] _next_pc_T_33 = io_now_pc + _GEN_6214; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [31:0] _next_pc_T_34 = io_now_pc + _GEN_6214; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [31:0] _GEN_6024 = ~global_data_setpc ? _next_pc_T_34 : _GEN_4943; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 150:30 154:17]
  wire [31:0] _event_exceptionInst_T = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _mstatusOld_WIRE_5 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusOld_2_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [7:0] mstatusOld_2_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [31:0] _mstatusNew_WIRE_5 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusNew_2_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_43 = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_45 = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_47 = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_49 = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_50 = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] mstatusNew_2_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_52 = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] mstatusNew_2_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] mstatusNew_2_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [7:0] mstatusNew_2_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [30:0] _next_csr_scause_T = {26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_scause_T_1 = {1'h0,26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 252:29]
  wire  _GEN_6044 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 164:35 257:35]
  wire  _mstatusNew_WIRE_4_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_sie = delegS ? 1'h0 : mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_6073 = mstatusNew_2_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _mstatusNew_WIRE_4_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_42 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] next_csr_mstatus_lo_lo_lo_2 = {mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_46 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_WIRE_4_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _GEN_6064 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 174:35 189:35]
  wire  mstatusNew_2_mie = delegS & mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_6083 = mstatusNew_2_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_2 = {mstatusOld_pad2,mstatusNew_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_44 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [2:0] next_csr_mstatus_lo_lo_hi_2 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [4:0] next_csr_mstatus_lo_lo_2 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_48 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusOld_WIRE_4_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_43 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _GEN_6043 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusNew_WIRE_4_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_spie = delegS ? mstatusOld_sie : mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_6072 = mstatusNew_2_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] next_csr_mstatus_lo_hi_lo_2 = {mstatusOld_ube,mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _mstatusNew_WIRE_4_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_51 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _GEN_6042 = io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 162:35 255:35]
  wire  _mstatusNew_WIRE_4_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _GEN_6071 = delegS ? io_now_internal_privilegeMode : {{1'd0}, mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_spp = _GEN_6071[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:30]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_2 = {mstatusOld_vs,mstatusNew_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusOld_WIRE_4_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_45 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _GEN_6063 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusNew_2_mpie = delegS ? mstatusOld_mpie : mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_6082 = mstatusNew_2_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [3:0] next_csr_mstatus_lo_hi_hi_2 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [5:0] next_csr_mstatus_lo_hi_2 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,
    mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [10:0] next_csr_mstatus_lo_2 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,mstatusNew_2_spie
    ,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _mstatusNew_WIRE_4_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_53 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_WIRE_4_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _GEN_6062 = io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 172:35 187:35]
  wire [1:0] mstatusNew_2_mpp = delegS ? mstatusOld_mpp : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] _GEN_6081 = mstatusNew_2_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [3:0] next_csr_mstatus_hi_lo_lo_2 = {mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_56 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_WIRE_4_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_55 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_2 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _mstatusNew_WIRE_4_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_54 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [3:0] next_csr_mstatus_hi_lo_hi_2 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [7:0] next_csr_mstatus_hi_lo_2 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_59 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_WIRE_4_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_58 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_2 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_57 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [2:0] next_csr_mstatus_hi_hi_lo_2 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_62 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [7:0] _mstatusNew_WIRE_4_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [7:0] _mstatusNew_T_61 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_2 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_60 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [9:0] next_csr_mstatus_hi_hi_hi_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [12:0] next_csr_mstatus_hi_hi_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [20:0] next_csr_mstatus_hi_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [31:0] _next_csr_mstatus_T_38 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _T_1124 = 5'h2 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [1:0] _T_1125 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:20]
  wire  _T_1126 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:27]
  wire [15:0] _next_csr_stval_T = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:69]
  wire [31:0] _next_csr_stval_T_1 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_6027 = inst[1:0] != 2'h3 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:{45,62} 272:41]
  wire  _T_1127 = 5'h1 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [1:0] _T_1128 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:20]
  wire  _T_1129 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:27]
  wire [15:0] _next_csr_stval_T_2 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:69]
  wire [31:0] _next_csr_stval_T_3 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_6028 = _T_1126 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:{45,62} 276:41]
  wire  _T_1130 = 5'h3 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [1:0] _T_1131 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:20]
  wire  _T_1132 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:27]
  wire [15:0] _next_csr_stval_T_4 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:69]
  wire [31:0] _next_csr_stval_T_5 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_6029 = _T_1126 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:{45,62} 281:41]
  wire  _T_1133 = 5'hb == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire  _T_1134 = 5'h6 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire  _T_1135 = 5'h4 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire  _T_1136 = 5'h0 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] mem_read_addr = io_valid ? _GEN_2708 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_6159 = mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_6030 = 5'h4 == exceptionNO ? mem_read_addr : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 296:26 259:35]
  wire [31:0] mem_write_addr = io_valid ? _GEN_2815 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_6166 = mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_6031 = 5'h6 == exceptionNO ? mem_write_addr : _GEN_6030; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 292:26]
  wire [31:0] _GEN_6032 = 5'hb == exceptionNO ? 32'h0 : _GEN_6031; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 288:26]
  wire [31:0] _GEN_6033 = 5'h3 == exceptionNO ? _GEN_6027 : _GEN_6032; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] _GEN_6034 = 5'h1 == exceptionNO ? _GEN_6027 : _GEN_6033; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] _GEN_6035 = 5'h2 == exceptionNO ? _GEN_6027 : _GEN_6034; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [29:0] _next_pc_T_35 = io_now_csr_stvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:46]
  wire [31:0] _next_pc_T_36 = {io_now_csr_stvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:62]
  wire [29:0] _next_pc_T_37 = io_now_csr_stvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:45]
  wire [31:0] _next_pc_T_38 = {27'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_6215 = {{2'd0}, io_now_csr_stvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [32:0] _next_pc_T_39 = _GEN_6215 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [31:0] _next_pc_T_40 = _GEN_6215 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [33:0] _next_pc_T_41 = {_next_pc_T_40, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:92]
  wire [33:0] _GEN_6037 = 2'h1 == io_now_csr_stvec[1:0] ? _next_pc_T_41 : {{2'd0}, _GEN_6024}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 317:29]
  wire [33:0] _GEN_6039 = 2'h0 == io_now_csr_stvec[1:0] ? {{2'd0}, _next_pc_T_36} : _GEN_6037; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 312:29]
  wire  _T_1140 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] now_csr_scause = io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6040 = 8'h20 == io_now_csr_MXLEN ? _next_csr_scause_T_1 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 252:23]
  wire  _GEN_6045 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 165:35 258:35]
  wire [31:0] now_csr_stval = io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6046 = 8'h20 == io_now_csr_MXLEN ? _GEN_6035 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] _GEN_6047 = 8'h20 == io_now_csr_MXLEN ? _next_csr_mstatus_T_38 : _GEN_6015; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 260:35]
  wire [33:0] _GEN_6049 = 8'h20 == io_now_csr_MXLEN ? _GEN_6039 : {{2'd0}, _GEN_6024}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [30:0] _next_csr_mcause_T_36 = {26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mcause_T_37 = {1'h0,26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 185:41]
  wire [1:0] next_csr_mstatus_lo_lo_lo_3 = {mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_3 = {mstatusOld_pad2,mstatusNew_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [2:0] next_csr_mstatus_lo_lo_hi_3 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [4:0] next_csr_mstatus_lo_lo_3 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_lo_hi_lo_3 = {mstatusOld_ube,mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_3 = {mstatusOld_vs,mstatusNew_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [3:0] next_csr_mstatus_lo_hi_hi_3 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [5:0] next_csr_mstatus_lo_hi_3 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,
    mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [10:0] next_csr_mstatus_lo_3 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,mstatusNew_2_spie
    ,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [3:0] next_csr_mstatus_hi_lo_lo_3 = {mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_3 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [3:0] next_csr_mstatus_hi_lo_hi_3 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [7:0] next_csr_mstatus_hi_lo_3 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_3 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [2:0] next_csr_mstatus_hi_hi_lo_3 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_3 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [9:0] next_csr_mstatus_hi_hi_hi_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [12:0] next_csr_mstatus_hi_hi_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [20:0] next_csr_mstatus_hi_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [31:0] _next_csr_mstatus_T_39 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire  _T_1142 = 5'h2 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1143 = 5'h1 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [1:0] _T_1144 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:20]
  wire  _T_1145 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:27]
  wire [15:0] _next_csr_mtval_T_54 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:69]
  wire [31:0] _next_csr_mtval_T_55 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_6050 = _T_1126 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:{45,62} 205:41]
  wire  _T_1146 = 5'hb == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1147 = 5'h6 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1148 = 5'h4 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1149 = 5'h0 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1150 = 5'h7 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1151 = 5'hd == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_1152 = 5'hc == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [31:0] _GEN_6051 = _T_1135 ? mem_read_addr : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 192:24 196:29 215:26]
  wire [31:0] _GEN_6052 = _T_1134 ? mem_write_addr : _GEN_6030; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 211:26]
  wire [31:0] _GEN_6053 = _T_1133 ? 32'h0 : _GEN_6031; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 208:26]
  wire [31:0] _GEN_6054 = _T_1127 ? _GEN_6027 : _GEN_6032; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [31:0] _GEN_6055 = _T_1124 ? 32'h0 : _GEN_6054; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 199:26]
  wire [29:0] _next_pc_T_42 = io_now_csr_mtvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:46]
  wire [31:0] _next_pc_T_43 = {io_now_csr_mtvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:62]
  wire [29:0] _next_pc_T_44 = io_now_csr_mtvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:45]
  wire [31:0] _next_pc_T_45 = {27'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_6216 = {{2'd0}, io_now_csr_mtvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [32:0] _next_pc_T_46 = _GEN_6216 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [31:0] _next_pc_T_47 = _GEN_6216 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [33:0] _next_pc_T_48 = {_next_pc_T_47, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:92]
  wire [33:0] _GEN_6057 = 2'h1 == io_now_csr_mtvec[1:0] ? _next_pc_T_48 : {{2'd0}, _GEN_6024}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 243:29]
  wire [33:0] _GEN_6059 = 2'h0 == io_now_csr_mtvec[1:0] ? {{2'd0}, _next_pc_T_43} : _GEN_6057; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 238:29]
  wire  _T_1156 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_6060 = _T_1123 ? _next_csr_scause_T_1 : _GEN_6022; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 185:35]
  wire [1:0] _GEN_6065 = 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 175:35 190:35]
  wire [31:0] _GEN_6066 = _T_1123 ? _GEN_6055 : _GEN_6023; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_6067 = _T_1123 ? _next_csr_mstatus_T_38 : _GEN_6015; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 193:24]
  wire [33:0] _GEN_6069 = _T_1123 ? _GEN_6059 : {{2'd0}, _GEN_6024}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_6075 = delegS ? _GEN_6040 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_6092 = raiseExceptionIntr ? _GEN_6075 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_scause = io_valid ? _GEN_6092 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6204 = next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6084 = delegS ? _GEN_6022 : _GEN_6060; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [31:0] _GEN_6098 = raiseExceptionIntr ? _GEN_6084 : _GEN_6022; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_mcause = io_valid ? _GEN_6098 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6199 = next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6070 = delegS ? next_csr_scause : next_csr_mcause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 161:35 171:35]
  wire [1:0] _GEN_6074 = delegS ? 2'h1 : 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [31:0] _GEN_6077 = delegS ? _GEN_6046 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_6078 = delegS ? _GEN_6047 : _GEN_6047; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [33:0] _GEN_6080 = delegS ? _GEN_6049 : _GEN_6069; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [31:0] _GEN_6086 = delegS ? _GEN_6023 : _GEN_6066; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [1:0] next_csr_mstatus_lo_lo_lo_4 = {mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_4 = {mstatusOld_pad2,mstatusNew_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [2:0] next_csr_mstatus_lo_lo_hi_4 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [4:0] next_csr_mstatus_lo_lo_4 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_lo_hi_lo_4 = {mstatusOld_ube,mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_4 = {mstatusOld_vs,mstatusNew_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [3:0] next_csr_mstatus_lo_hi_hi_4 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [5:0] next_csr_mstatus_lo_hi_4 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,
    mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [10:0] next_csr_mstatus_lo_4 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,mstatusNew_2_spie
    ,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [3:0] next_csr_mstatus_hi_lo_lo_4 = {mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_4 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [3:0] next_csr_mstatus_hi_lo_hi_4 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [7:0] next_csr_mstatus_hi_lo_4 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_4 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [2:0] next_csr_mstatus_hi_hi_lo_4 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_4 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [9:0] next_csr_mstatus_hi_hi_hi_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [12:0] next_csr_mstatus_hi_hi_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [20:0] next_csr_mstatus_hi_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [31:0] _next_csr_mstatus_T_40 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire  _GEN_6087 = raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [31:0] _event_WIRE_cause = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_6088 = raiseExceptionIntr ? _GEN_6070 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _event_WIRE_exceptionPC = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_6089 = raiseExceptionIntr ? io_now_pc : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 151:25]
  wire [31:0] _event_WIRE_exceptionInst = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_6090 = raiseExceptionIntr ? inst : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 152:25]
  wire [1:0] _GEN_6091 = raiseExceptionIntr ? _GEN_6074 : _GEN_4939; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _GEN_6094 = raiseExceptionIntr ? _GEN_6077 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _GEN_6095 = raiseExceptionIntr ? _next_csr_mstatus_T_38 : _GEN_6015; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 181:22]
  wire [33:0] _GEN_6097 = raiseExceptionIntr ? _GEN_6080 : {{2'd0}, _GEN_6024}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _GEN_6100 = raiseExceptionIntr ? _GEN_6086 : _GEN_6023; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_cycle = io_valid ? _next_csr_cycle_T_1 : io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 126:20 111:21]
  wire [31:0] _GEN_6104 = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 131:16 115:21]
  wire [2:0] funct3 = io_valid ? _GEN_5975 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 18:24]
  wire [6:0] opcode = io_valid ? _GEN_5977 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 16:24]
  wire [31:0] next_reg_0 = io_valid ? 32'h0 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  wire [31:0] next_reg_1 = io_valid ? _GEN_5983 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_2 = io_valid ? _GEN_5984 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_3 = io_valid ? _GEN_5985 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_4 = io_valid ? _GEN_5986 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_5 = io_valid ? _GEN_5987 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_6 = io_valid ? _GEN_5988 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_7 = io_valid ? _GEN_5989 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_8 = io_valid ? _GEN_5990 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_9 = io_valid ? _GEN_5991 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_10 = io_valid ? _GEN_5992 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_11 = io_valid ? _GEN_5993 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_12 = io_valid ? _GEN_5994 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_13 = io_valid ? _GEN_5995 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_14 = io_valid ? _GEN_5996 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_15 = io_valid ? _GEN_5997 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_16 = io_valid ? _GEN_5998 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_17 = io_valid ? _GEN_5999 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_18 = io_valid ? _GEN_6000 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_19 = io_valid ? _GEN_6001 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_20 = io_valid ? _GEN_6002 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_21 = io_valid ? _GEN_6003 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_22 = io_valid ? _GEN_6004 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_23 = io_valid ? _GEN_6005 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_24 = io_valid ? _GEN_6006 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_25 = io_valid ? _GEN_6007 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_26 = io_valid ? _GEN_6008 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_27 = io_valid ? _GEN_6009 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_28 = io_valid ? _GEN_6010 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_29 = io_valid ? _GEN_6011 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_30 = io_valid ? _GEN_6012 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_31 = io_valid ? _GEN_6013 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [6:0] funct7 = io_valid ? _GEN_4862 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 21:24]
  wire [33:0] _GEN_6151 = io_valid ? _GEN_6097 : {{2'd0}, io_now_pc}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mtval = io_valid ? _GEN_6100 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  mem_read_valid = io_valid & _GEN_2707; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] mem_read_memWidth = io_valid ? _GEN_2709 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  mem_write_valid = io_valid & _GEN_2814; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] mem_write_memWidth = io_valid ? _GEN_2816 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] mem_write_data = io_valid ? _GEN_2817 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  ph1 = io_valid & _GEN_4327; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:22]
  wire [4:0] ph5 = io_valid ? _GEN_4329 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:52]
  wire [1:0] op = io_valid ? _GEN_4330 : 2'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 97:24]
  wire [5:0] ph6 = io_valid ? _GEN_2627 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 104:22]
  wire [2:0] ph3 = io_valid ? _GEN_3607 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:22]
  wire [1:0] ph2 = io_valid ? _GEN_2810 : 2'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:52]
  wire [10:0] ph11 = io_valid ? _GEN_2827 : 11'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 107:22]
  wire [3:0] funct4 = io_valid ? _GEN_3748 : 4'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 95:24]
  wire [7:0] ph8 = io_valid ? _GEN_3226 : 8'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 105:22]
  wire [5:0] funct6 = io_valid ? _GEN_4287 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 96:24]
  wire [1:0] funct2 = io_valid ? _GEN_4289 : 2'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 94:24]
  wire [1:0] next_internal_privilegeMode = io_valid ? _GEN_6091 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mstatus = io_valid ? _GEN_6095 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6190 = retTarget; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] next_csr_misa = io_valid ? _GEN_6014 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mscratch = io_valid ? _GEN_6016 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mtvec = io_valid ? _GEN_6017 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mcounteren = io_valid ? _GEN_6018 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mip = io_valid ? _GEN_6019 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mie = io_valid ? _GEN_6020 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  _event_WIRE_valid = 1'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire  event_valid = io_valid & raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] event_cause = io_valid ? _GEN_6088 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] event_exceptionPC = io_valid ? _GEN_6089 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] event_exceptionInst = io_valid ? _GEN_6090 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] next_csr_stval = io_valid ? _GEN_6094 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] now_csr_mstatush = io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mideleg = io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_scounteren = io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_sscratch = io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg0 = io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg1 = io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg2 = io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg3 = io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr0 = io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr1 = io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr2 = io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr3 = io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] now_csr_ILEN = io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6111 = next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  wire [31:0] _GEN_6112 = next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6113 = next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6114 = next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6115 = next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6116 = next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6117 = next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6118 = next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6119 = next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6120 = next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6121 = next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6122 = next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6123 = next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6124 = next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6125 = next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6126 = next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6127 = next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6128 = next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6129 = next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6130 = next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6131 = next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6132 = next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6133 = next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6134 = next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6135 = next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6136 = next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6137 = next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6138 = next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6139 = next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6140 = next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6141 = next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6142 = next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_pc = _GEN_6151[31:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 18:18]
  wire [31:0] _GEN_6192 = next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6189 = next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mstatush = io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6193 = next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6194 = next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6195 = next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mideleg = io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6196 = next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6197 = next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6152 = next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_6101 = next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 126:20 111:21]
  wire [31:0] next_csr_scounteren = io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_6206 = next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_sscratch = io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg0 = io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg1 = io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg2 = io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg3 = io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr0 = io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr1 = io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr2 = io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr3 = io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] next_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] next_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] next_csr_ILEN = io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [1:0] _GEN_6188 = next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] iFetchpc = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 131:16 115:21]
  wire  _GEN_6158 = mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] _GEN_6160 = mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  _GEN_6165 = mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] _GEN_6167 = mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_6168 = mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  _GEN_6200 = event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] _event_WIRE_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] event_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_6201 = event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] _GEN_6202 = event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] _GEN_6203 = event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire  _exceptionVec_WIRE_10 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _exceptionVec_WIRE_14 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_10 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_14 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [6:0] _GEN_6109 = opcode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 16:24]
  wire [2:0] _GEN_6107 = funct3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 18:24]
  wire [6:0] _GEN_6144 = funct7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 21:24]
  wire [1:0] _GEN_6186 = funct2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 94:24]
  wire [3:0] _GEN_6183 = funct4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 95:24]
  wire [5:0] _GEN_6185 = funct6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 96:24]
  wire [1:0] _GEN_6175 = op; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 97:24]
  wire  _GEN_6173 = ph1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:22]
  wire [4:0] _GEN_6174 = ph5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:52]
  wire [5:0] _GEN_6176 = ph6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 104:22]
  wire [7:0] _GEN_6184 = ph8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 105:22]
  wire [2:0] _GEN_6177 = ph3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:22]
  wire [1:0] _GEN_6179 = ph2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:52]
  wire [10:0] _GEN_6182 = ph11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 107:22]
  wire [31:0] _GEN_4941 = retTarget; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _mem_WIRE_read_data = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire  _mstatusOld_WIRE_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [7:0] _mstatusOld_WIRE_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_20 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [7:0] _mstatusOld_T_19 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_17 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_16 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_15 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_14 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_13 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_12 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_11 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_10 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_9 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_7 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_6 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_4 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_3 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_2 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_1 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_2_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [7:0] _mstatusOld_WIRE_2_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_WIRE_2_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_WIRE_2_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_WIRE_2_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_41 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [7:0] _mstatusOld_T_40 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_39 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_38 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_37 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_36 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_35 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_34 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_33 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_32 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_30 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_29 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_27 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_26 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_25 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_24 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_23 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_22 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_21 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusNew_WIRE_2_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusOld_WIRE_4_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [7:0] _mstatusOld_WIRE_4_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_62 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [7:0] _mstatusOld_T_61 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_60 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_59 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_58 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_57 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_56 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_55 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_54 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_53 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_52 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_51 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_50 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_49 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_48 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_47 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_46 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_44 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_42 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  assign io_iFetchpc = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 131:16 115:21]
  assign io_mem_read_valid = io_valid & _GEN_2707; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_addr = io_valid ? _GEN_2708 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_memWidth = io_valid ? _GEN_2709 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_valid = io_valid & _GEN_2814; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_addr = io_valid ? _GEN_2815 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_memWidth = io_valid ? _GEN_2816 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_data = io_valid ? _GEN_2817 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_next_reg_0 = io_valid ? 32'h0 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  assign io_next_reg_1 = io_valid ? _GEN_5983 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_2 = io_valid ? _GEN_5984 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_3 = io_valid ? _GEN_5985 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_4 = io_valid ? _GEN_5986 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_5 = io_valid ? _GEN_5987 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_6 = io_valid ? _GEN_5988 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_7 = io_valid ? _GEN_5989 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_8 = io_valid ? _GEN_5990 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_9 = io_valid ? _GEN_5991 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_10 = io_valid ? _GEN_5992 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_11 = io_valid ? _GEN_5993 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_12 = io_valid ? _GEN_5994 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_13 = io_valid ? _GEN_5995 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_14 = io_valid ? _GEN_5996 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_15 = io_valid ? _GEN_5997 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_16 = io_valid ? _GEN_5998 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_17 = io_valid ? _GEN_5999 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_18 = io_valid ? _GEN_6000 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_19 = io_valid ? _GEN_6001 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_20 = io_valid ? _GEN_6002 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_21 = io_valid ? _GEN_6003 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_22 = io_valid ? _GEN_6004 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_23 = io_valid ? _GEN_6005 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_24 = io_valid ? _GEN_6006 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_25 = io_valid ? _GEN_6007 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_26 = io_valid ? _GEN_6008 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_27 = io_valid ? _GEN_6009 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_28 = io_valid ? _GEN_6010 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_29 = io_valid ? _GEN_6011 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_30 = io_valid ? _GEN_6012 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_31 = io_valid ? _GEN_6013 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_pc = _GEN_6151[31:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 18:18]
  assign io_next_csr_misa = io_valid ? _GEN_6014 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mstatus = io_valid ? _GEN_6095 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mstatush = io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mscratch = io_valid ? _GEN_6016 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mtvec = io_valid ? _GEN_6017 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mcounteren = io_valid ? _GEN_6018 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mideleg = io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mip = io_valid ? _GEN_6019 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mie = io_valid ? _GEN_6020 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mepc = io_valid ? _GEN_6099 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mcause = io_valid ? _GEN_6098 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mtval = io_valid ? _GEN_6100 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_cycle = io_valid ? _next_csr_cycle_T_1 : io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 126:20 111:21]
  assign io_next_csr_scounteren = io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_scause = io_valid ? _GEN_6092 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_sepc = io_valid ? _GEN_6093 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_stval = io_valid ? _GEN_6094 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_sscratch = io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg0 = io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg1 = io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg2 = io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg3 = io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr0 = io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr1 = io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr2 = io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr3 = io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_ILEN = io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_internal_privilegeMode = io_valid ? _GEN_6091 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_event_valid = io_valid & raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  assign io_event_cause = io_valid ? _GEN_6088 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionPC = io_valid ? _GEN_6089 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionInst = io_valid ? _GEN_6090 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
endmodule
module RiscvCore(
  input         clock,
  input         reset,
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_iFetchpc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_now_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_now_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_now_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [1:0]  io_now_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_next_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_next_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_next_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [1:0]  io_next_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
`endif // RANDOMIZE_REG_INIT
  wire  trans_clock; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_reset; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_iFetchpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [5:0] trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [5:0] trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_intrNO; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [30:0] _state_state_csr_misaInitVal_T = 31'h40000000; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 335:25]
  wire  _state_state_csr_misaInitVal_T_1 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire  _state_state_csr_misaInitVal_T_2 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [8:0] _state_state_csr_misaInitVal_T_3 = 9'h100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire [8:0] _state_state_csr_misaInitVal_T_4 = 9'h101; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [12:0] _state_state_csr_misaInitVal_T_5 = 13'h1000; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire [12:0] _state_state_csr_misaInitVal_T_6 = 13'h1101; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [2:0] _state_state_csr_misaInitVal_T_7 = 3'h4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire [12:0] _state_state_csr_misaInitVal_T_8 = 13'h1105; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [20:0] _state_state_csr_misaInitVal_T_9 = 21'h100000; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire [20:0] _state_state_csr_misaInitVal_T_10 = 21'h101105; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [30:0] state_state_csr_misaInitVal = 31'h40101105; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:20]
  wire [31:0] state_state_csr_csr_mstatus = 32'h1800; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 353:17]
  wire [31:0] _state_state_csr_mstatusStruct_WIRE = 32'h1800; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 353:17]
  wire  _state_state_csr_mstatusStruct_T = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_2 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_3 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_4 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_5 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_6 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_7 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_8 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_9 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_10 = 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_11 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_12 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_13 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_14 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_15 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_16 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_17 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_18 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [7:0] _state_state_csr_mstatusStruct_T_19 = 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_20 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  reg [31:0] state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [1:0] state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  wire [31:0] state_state_reg_0 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_1 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_2 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_3 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_4 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_5 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_6 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_7 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_8 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_9 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_10 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_11 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_12 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_13 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_14 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_15 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_16 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_17 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_18 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_19 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_20 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_21 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_22 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_23 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_24 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_25 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_26 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_27 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_28 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_29 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_30 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_31 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_pc = 32'h8000; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 84:15]
  wire [31:0] state_state_csr_csr_misa = 32'h40101105; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 343:14]
  wire [31:0] state_state_csr_misa = 32'h40101105; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 343:14]
  wire [31:0] state_state_csr_csr_mvendorid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 347:19]
  wire [31:0] state_state_csr_mvendorid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 347:19]
  wire [31:0] state_state_csr_csr_marchid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 349:17]
  wire [31:0] state_state_csr_marchid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 349:17]
  wire [31:0] state_state_csr_csr_mimpid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 351:17]
  wire [31:0] state_state_csr_mimpid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 351:17]
  wire [31:0] state_state_csr_csr_mhartid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 352:17]
  wire [31:0] state_state_csr_mhartid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 352:17]
  wire [31:0] state_state_csr_mstatus = 32'h1800; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 353:17]
  wire [31:0] state_state_csr_csr_mstatush = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 357:20]
  wire [31:0] state_state_csr_mstatush = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 357:20]
  wire [31:0] state_state_csr_csr_mscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 358:20]
  wire [31:0] state_state_csr_mscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 358:20]
  wire [31:0] state_state_csr_csr_mtvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 359:20]
  wire [31:0] state_state_csr_mtvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 359:20]
  wire [31:0] state_state_csr_csr_mcounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 360:20]
  wire [31:0] state_state_csr_mcounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 360:20]
  wire [31:0] state_state_csr_csr_medeleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 361:20]
  wire [31:0] state_state_csr_medeleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 361:20]
  wire [31:0] state_state_csr_csr_mideleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 362:20]
  wire [31:0] state_state_csr_mideleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 362:20]
  wire [31:0] state_state_csr_csr_mip = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 363:20]
  wire [31:0] state_state_csr_mip = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 363:20]
  wire [31:0] state_state_csr_csr_mie = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 364:20]
  wire [31:0] state_state_csr_mie = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 364:20]
  wire [31:0] state_state_csr_csr_mepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 365:20]
  wire [31:0] state_state_csr_mepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 365:20]
  wire [31:0] state_state_csr_csr_mcause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 366:20]
  wire [31:0] state_state_csr_mcause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 366:20]
  wire [31:0] state_state_csr_csr_mtval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 367:20]
  wire [31:0] state_state_csr_mtval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 367:20]
  wire [31:0] state_state_csr_csr_cycle = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 368:20]
  wire [31:0] state_state_csr_cycle = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 368:20]
  wire [31:0] state_state_csr_csr_scounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 372:20]
  wire [31:0] state_state_csr_scounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 372:20]
  wire [31:0] state_state_csr_csr_scause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 371:20]
  wire [31:0] state_state_csr_scause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 371:20]
  wire [31:0] state_state_csr_csr_stvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 373:20]
  wire [31:0] state_state_csr_stvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 373:20]
  wire [31:0] state_state_csr_csr_sepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 374:20]
  wire [31:0] state_state_csr_sepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 374:20]
  wire [31:0] state_state_csr_csr_stval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 375:20]
  wire [31:0] state_state_csr_stval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 375:20]
  wire [31:0] state_state_csr_csr_sscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 376:20]
  wire [31:0] state_state_csr_sscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 376:20]
  wire [31:0] state_state_csr_csr_satp = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 378:14]
  wire [31:0] state_state_csr_satp = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 378:14]
  wire [31:0] state_state_csr_csr_pmpcfg0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 386:18]
  wire [31:0] state_state_csr_pmpcfg0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 386:18]
  wire [31:0] state_state_csr_csr_pmpcfg1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 387:18]
  wire [31:0] state_state_csr_pmpcfg1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 387:18]
  wire [31:0] state_state_csr_csr_pmpcfg2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 388:18]
  wire [31:0] state_state_csr_pmpcfg2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 388:18]
  wire [31:0] state_state_csr_csr_pmpcfg3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 389:18]
  wire [31:0] state_state_csr_pmpcfg3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 389:18]
  wire [31:0] state_state_csr_csr_pmpaddr0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 390:18]
  wire [31:0] state_state_csr_pmpaddr0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 390:18]
  wire [31:0] state_state_csr_csr_pmpaddr1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 391:18]
  wire [31:0] state_state_csr_pmpaddr1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 391:18]
  wire [31:0] state_state_csr_csr_pmpaddr2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 392:18]
  wire [31:0] state_state_csr_pmpaddr2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 392:18]
  wire [31:0] state_state_csr_csr_pmpaddr3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 393:18]
  wire [31:0] state_state_csr_pmpaddr3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 393:18]
  wire [7:0] state_state_csr_csr_MXLEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 398:15]
  wire [7:0] state_state_csr_MXLEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 398:15]
  wire [7:0] state_state_csr_csr_IALIGN = 8'h10; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 399:16]
  wire [7:0] state_state_csr_IALIGN = 8'h10; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 399:16]
  wire [7:0] state_state_csr_csr_ILEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 403:14]
  wire [7:0] state_state_csr_ILEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 403:14]
  wire [1:0] state_state_internal_internal_privilegeMode = 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 61:24 62:28]
  wire [1:0] state_state_internal_privilegeMode = 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 61:24 62:28]
  wire  state_state_csr_mstatusStruct_sd = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [7:0] state_state_csr_mstatusStruct_pad0 = 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_tsr = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_tw = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_tvm = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mxr = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_sum = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mprv = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_xs = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_fs = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_mpp = 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_vs = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_spp = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mpie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_ube = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_spie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_pad2 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_pad3 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_sie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_pad4 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  RiscvTrans trans ( // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
    .clock(trans_clock),
    .reset(trans_reset),
    .io_inst(trans_io_inst),
    .io_valid(trans_io_valid),
    .io_iFetchpc(trans_io_iFetchpc),
    .io_mem_read_valid(trans_io_mem_read_valid),
    .io_mem_read_addr(trans_io_mem_read_addr),
    .io_mem_read_memWidth(trans_io_mem_read_memWidth),
    .io_mem_read_data(trans_io_mem_read_data),
    .io_mem_write_valid(trans_io_mem_write_valid),
    .io_mem_write_addr(trans_io_mem_write_addr),
    .io_mem_write_memWidth(trans_io_mem_write_memWidth),
    .io_mem_write_data(trans_io_mem_write_data),
    .io_now_reg_0(trans_io_now_reg_0),
    .io_now_reg_1(trans_io_now_reg_1),
    .io_now_reg_2(trans_io_now_reg_2),
    .io_now_reg_3(trans_io_now_reg_3),
    .io_now_reg_4(trans_io_now_reg_4),
    .io_now_reg_5(trans_io_now_reg_5),
    .io_now_reg_6(trans_io_now_reg_6),
    .io_now_reg_7(trans_io_now_reg_7),
    .io_now_reg_8(trans_io_now_reg_8),
    .io_now_reg_9(trans_io_now_reg_9),
    .io_now_reg_10(trans_io_now_reg_10),
    .io_now_reg_11(trans_io_now_reg_11),
    .io_now_reg_12(trans_io_now_reg_12),
    .io_now_reg_13(trans_io_now_reg_13),
    .io_now_reg_14(trans_io_now_reg_14),
    .io_now_reg_15(trans_io_now_reg_15),
    .io_now_reg_16(trans_io_now_reg_16),
    .io_now_reg_17(trans_io_now_reg_17),
    .io_now_reg_18(trans_io_now_reg_18),
    .io_now_reg_19(trans_io_now_reg_19),
    .io_now_reg_20(trans_io_now_reg_20),
    .io_now_reg_21(trans_io_now_reg_21),
    .io_now_reg_22(trans_io_now_reg_22),
    .io_now_reg_23(trans_io_now_reg_23),
    .io_now_reg_24(trans_io_now_reg_24),
    .io_now_reg_25(trans_io_now_reg_25),
    .io_now_reg_26(trans_io_now_reg_26),
    .io_now_reg_27(trans_io_now_reg_27),
    .io_now_reg_28(trans_io_now_reg_28),
    .io_now_reg_29(trans_io_now_reg_29),
    .io_now_reg_30(trans_io_now_reg_30),
    .io_now_reg_31(trans_io_now_reg_31),
    .io_now_pc(trans_io_now_pc),
    .io_now_csr_misa(trans_io_now_csr_misa),
    .io_now_csr_mvendorid(trans_io_now_csr_mvendorid),
    .io_now_csr_marchid(trans_io_now_csr_marchid),
    .io_now_csr_mimpid(trans_io_now_csr_mimpid),
    .io_now_csr_mhartid(trans_io_now_csr_mhartid),
    .io_now_csr_mstatus(trans_io_now_csr_mstatus),
    .io_now_csr_mstatush(trans_io_now_csr_mstatush),
    .io_now_csr_mscratch(trans_io_now_csr_mscratch),
    .io_now_csr_mtvec(trans_io_now_csr_mtvec),
    .io_now_csr_mcounteren(trans_io_now_csr_mcounteren),
    .io_now_csr_medeleg(trans_io_now_csr_medeleg),
    .io_now_csr_mideleg(trans_io_now_csr_mideleg),
    .io_now_csr_mip(trans_io_now_csr_mip),
    .io_now_csr_mie(trans_io_now_csr_mie),
    .io_now_csr_mepc(trans_io_now_csr_mepc),
    .io_now_csr_mcause(trans_io_now_csr_mcause),
    .io_now_csr_mtval(trans_io_now_csr_mtval),
    .io_now_csr_cycle(trans_io_now_csr_cycle),
    .io_now_csr_scounteren(trans_io_now_csr_scounteren),
    .io_now_csr_scause(trans_io_now_csr_scause),
    .io_now_csr_stvec(trans_io_now_csr_stvec),
    .io_now_csr_sepc(trans_io_now_csr_sepc),
    .io_now_csr_stval(trans_io_now_csr_stval),
    .io_now_csr_sscratch(trans_io_now_csr_sscratch),
    .io_now_csr_satp(trans_io_now_csr_satp),
    .io_now_csr_pmpcfg0(trans_io_now_csr_pmpcfg0),
    .io_now_csr_pmpcfg1(trans_io_now_csr_pmpcfg1),
    .io_now_csr_pmpcfg2(trans_io_now_csr_pmpcfg2),
    .io_now_csr_pmpcfg3(trans_io_now_csr_pmpcfg3),
    .io_now_csr_pmpaddr0(trans_io_now_csr_pmpaddr0),
    .io_now_csr_pmpaddr1(trans_io_now_csr_pmpaddr1),
    .io_now_csr_pmpaddr2(trans_io_now_csr_pmpaddr2),
    .io_now_csr_pmpaddr3(trans_io_now_csr_pmpaddr3),
    .io_now_csr_MXLEN(trans_io_now_csr_MXLEN),
    .io_now_csr_IALIGN(trans_io_now_csr_IALIGN),
    .io_now_csr_ILEN(trans_io_now_csr_ILEN),
    .io_now_internal_privilegeMode(trans_io_now_internal_privilegeMode),
    .io_next_reg_0(trans_io_next_reg_0),
    .io_next_reg_1(trans_io_next_reg_1),
    .io_next_reg_2(trans_io_next_reg_2),
    .io_next_reg_3(trans_io_next_reg_3),
    .io_next_reg_4(trans_io_next_reg_4),
    .io_next_reg_5(trans_io_next_reg_5),
    .io_next_reg_6(trans_io_next_reg_6),
    .io_next_reg_7(trans_io_next_reg_7),
    .io_next_reg_8(trans_io_next_reg_8),
    .io_next_reg_9(trans_io_next_reg_9),
    .io_next_reg_10(trans_io_next_reg_10),
    .io_next_reg_11(trans_io_next_reg_11),
    .io_next_reg_12(trans_io_next_reg_12),
    .io_next_reg_13(trans_io_next_reg_13),
    .io_next_reg_14(trans_io_next_reg_14),
    .io_next_reg_15(trans_io_next_reg_15),
    .io_next_reg_16(trans_io_next_reg_16),
    .io_next_reg_17(trans_io_next_reg_17),
    .io_next_reg_18(trans_io_next_reg_18),
    .io_next_reg_19(trans_io_next_reg_19),
    .io_next_reg_20(trans_io_next_reg_20),
    .io_next_reg_21(trans_io_next_reg_21),
    .io_next_reg_22(trans_io_next_reg_22),
    .io_next_reg_23(trans_io_next_reg_23),
    .io_next_reg_24(trans_io_next_reg_24),
    .io_next_reg_25(trans_io_next_reg_25),
    .io_next_reg_26(trans_io_next_reg_26),
    .io_next_reg_27(trans_io_next_reg_27),
    .io_next_reg_28(trans_io_next_reg_28),
    .io_next_reg_29(trans_io_next_reg_29),
    .io_next_reg_30(trans_io_next_reg_30),
    .io_next_reg_31(trans_io_next_reg_31),
    .io_next_pc(trans_io_next_pc),
    .io_next_csr_misa(trans_io_next_csr_misa),
    .io_next_csr_mvendorid(trans_io_next_csr_mvendorid),
    .io_next_csr_marchid(trans_io_next_csr_marchid),
    .io_next_csr_mimpid(trans_io_next_csr_mimpid),
    .io_next_csr_mhartid(trans_io_next_csr_mhartid),
    .io_next_csr_mstatus(trans_io_next_csr_mstatus),
    .io_next_csr_mstatush(trans_io_next_csr_mstatush),
    .io_next_csr_mscratch(trans_io_next_csr_mscratch),
    .io_next_csr_mtvec(trans_io_next_csr_mtvec),
    .io_next_csr_mcounteren(trans_io_next_csr_mcounteren),
    .io_next_csr_medeleg(trans_io_next_csr_medeleg),
    .io_next_csr_mideleg(trans_io_next_csr_mideleg),
    .io_next_csr_mip(trans_io_next_csr_mip),
    .io_next_csr_mie(trans_io_next_csr_mie),
    .io_next_csr_mepc(trans_io_next_csr_mepc),
    .io_next_csr_mcause(trans_io_next_csr_mcause),
    .io_next_csr_mtval(trans_io_next_csr_mtval),
    .io_next_csr_cycle(trans_io_next_csr_cycle),
    .io_next_csr_scounteren(trans_io_next_csr_scounteren),
    .io_next_csr_scause(trans_io_next_csr_scause),
    .io_next_csr_stvec(trans_io_next_csr_stvec),
    .io_next_csr_sepc(trans_io_next_csr_sepc),
    .io_next_csr_stval(trans_io_next_csr_stval),
    .io_next_csr_sscratch(trans_io_next_csr_sscratch),
    .io_next_csr_satp(trans_io_next_csr_satp),
    .io_next_csr_pmpcfg0(trans_io_next_csr_pmpcfg0),
    .io_next_csr_pmpcfg1(trans_io_next_csr_pmpcfg1),
    .io_next_csr_pmpcfg2(trans_io_next_csr_pmpcfg2),
    .io_next_csr_pmpcfg3(trans_io_next_csr_pmpcfg3),
    .io_next_csr_pmpaddr0(trans_io_next_csr_pmpaddr0),
    .io_next_csr_pmpaddr1(trans_io_next_csr_pmpaddr1),
    .io_next_csr_pmpaddr2(trans_io_next_csr_pmpaddr2),
    .io_next_csr_pmpaddr3(trans_io_next_csr_pmpaddr3),
    .io_next_csr_MXLEN(trans_io_next_csr_MXLEN),
    .io_next_csr_IALIGN(trans_io_next_csr_IALIGN),
    .io_next_csr_ILEN(trans_io_next_csr_ILEN),
    .io_next_internal_privilegeMode(trans_io_next_internal_privilegeMode),
    .io_event_valid(trans_io_event_valid),
    .io_event_intrNO(trans_io_event_intrNO),
    .io_event_cause(trans_io_event_cause),
    .io_event_exceptionPC(trans_io_event_exceptionPC),
    .io_event_exceptionInst(trans_io_event_exceptionInst)
  );
  assign io_iFetchpc = trans_io_iFetchpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 203:15]
  assign io_mem_read_valid = trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_addr = trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_memWidth = trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_valid = trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_addr = trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_memWidth = trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_data = trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_now_reg_0 = state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_1 = state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_2 = state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_3 = state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_4 = state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_5 = state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_6 = state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_7 = state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_8 = state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_9 = state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_10 = state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_11 = state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_12 = state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_13 = state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_14 = state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_15 = state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_16 = state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_17 = state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_18 = state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_19 = state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_20 = state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_21 = state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_22 = state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_23 = state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_24 = state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_25 = state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_26 = state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_27 = state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_28 = state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_29 = state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_30 = state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_31 = state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_misa = state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mvendorid = state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_marchid = state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mimpid = state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mhartid = state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mstatus = state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mstatush = state_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mscratch = state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mtvec = state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mcounteren = state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_medeleg = state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mideleg = state_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mip = state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mie = state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mepc = state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mcause = state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mtval = state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_cycle = state_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_scounteren = state_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_scause = state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_stvec = state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_sepc = state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_stval = state_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_sscratch = state_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_satp = state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg0 = state_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg1 = state_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg2 = state_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg3 = state_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr0 = state_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr1 = state_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr2 = state_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr3 = state_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_MXLEN = state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_IALIGN = state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_ILEN = state_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_internal_privilegeMode = state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_next_reg_0 = trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_1 = trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_2 = trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_3 = trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_4 = trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_5 = trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_6 = trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_7 = trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_8 = trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_9 = trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_10 = trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_11 = trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_12 = trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_13 = trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_14 = trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_15 = trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_16 = trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_17 = trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_18 = trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_19 = trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_20 = trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_21 = trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_22 = trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_23 = trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_24 = trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_25 = trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_26 = trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_27 = trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_28 = trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_29 = trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_30 = trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_31 = trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_pc = trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_misa = trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mvendorid = trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_marchid = trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mimpid = trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mhartid = trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mstatus = trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mstatush = trans_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mscratch = trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtvec = trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcounteren = trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_medeleg = trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mideleg = trans_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mip = trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mie = trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mepc = trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcause = trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtval = trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_cycle = trans_io_next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_scounteren = trans_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_scause = trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_stvec = trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_sepc = trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_stval = trans_io_next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_sscratch = trans_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_satp = trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg0 = trans_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg1 = trans_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg2 = trans_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg3 = trans_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr0 = trans_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr1 = trans_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr2 = trans_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr3 = trans_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_MXLEN = trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_IALIGN = trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_ILEN = trans_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_internal_privilegeMode = trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_event_valid = trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_cause = trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionPC = trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionInst = trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign trans_clock = clock;
  assign trans_reset = reset;
  assign trans_io_inst = io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 192:18]
  assign trans_io_valid = io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 193:18]
  assign trans_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign trans_io_now_reg_0 = state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_1 = state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_2 = state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_3 = state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_4 = state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_5 = state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_6 = state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_7 = state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_8 = state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_9 = state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_10 = state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_11 = state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_12 = state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_13 = state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_14 = state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_15 = state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_16 = state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_17 = state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_18 = state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_19 = state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_20 = state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_21 = state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_22 = state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_23 = state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_24 = state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_25 = state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_26 = state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_27 = state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_28 = state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_29 = state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_30 = state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_31 = state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_misa = state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mvendorid = state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_marchid = state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mimpid = state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mhartid = state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mstatus = state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mstatush = state_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mscratch = state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtvec = state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcounteren = state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_medeleg = state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mideleg = state_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mip = state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mie = state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mepc = state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcause = state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtval = state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_cycle = state_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_scounteren = state_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_scause = state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_stvec = state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_sepc = state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_stval = state_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_sscratch = state_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_satp = state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg0 = state_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg1 = state_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg2 = state_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg3 = state_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr0 = state_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr1 = state_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr2 = state_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr3 = state_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_MXLEN = state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_IALIGN = state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_ILEN = state_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_internal_privilegeMode = state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_0 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_0 <= trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_1 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_1 <= trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_2 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_2 <= trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_3 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_3 <= trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_4 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_4 <= trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_5 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_5 <= trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_6 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_6 <= trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_7 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_7 <= trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_8 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_8 <= trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_9 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_9 <= trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_10 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_10 <= trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_11 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_11 <= trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_12 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_12 <= trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_13 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_13 <= trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_14 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_14 <= trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_15 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_15 <= trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_16 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_16 <= trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_17 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_17 <= trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_18 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_18 <= trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_19 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_19 <= trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_20 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_20 <= trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_21 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_21 <= trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_22 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_22 <= trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_23 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_23 <= trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_24 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_24 <= trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_25 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_25 <= trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_26 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_26 <= trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_27 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_27 <= trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_28 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_28 <= trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_29 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_29 <= trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_30 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_30 <= trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_31 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_31 <= trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_pc <= 32'h8000; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_pc <= trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_misa <= 32'h40101105; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_misa <= trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mvendorid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mvendorid <= trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_marchid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_marchid <= trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mimpid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mimpid <= trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mhartid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mhartid <= trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mstatus <= 32'h1800; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mstatus <= trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mstatush <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mstatush <= trans_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mscratch <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mscratch <= trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtvec <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtvec <= trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcounteren <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcounteren <= trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_medeleg <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_medeleg <= trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mideleg <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mideleg <= trans_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mip <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mip <= trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mie <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mie <= trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mepc <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mepc <= trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcause <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcause <= trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtval <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtval <= trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_cycle <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_cycle <= trans_io_next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_scounteren <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_scounteren <= trans_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_scause <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_scause <= trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_stvec <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_stvec <= trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_sepc <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_sepc <= trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_stval <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_stval <= trans_io_next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_sscratch <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_sscratch <= trans_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_satp <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_satp <= trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg0 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg0 <= trans_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg1 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg1 <= trans_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg2 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg2 <= trans_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg3 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg3 <= trans_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr0 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr0 <= trans_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr1 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr1 <= trans_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr2 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr2 <= trans_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr3 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr3 <= trans_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_MXLEN <= 8'h20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_MXLEN <= trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_IALIGN <= 8'h10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_IALIGN <= trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_ILEN <= 8'h20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_ILEN <= trans_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_internal_privilegeMode <= 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_internal_privilegeMode <= trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  state_reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state_reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  state_reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  state_reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  state_reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  state_reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  state_reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  state_reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_reg_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  state_reg_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  state_reg_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  state_reg_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  state_reg_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  state_reg_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  state_reg_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  state_reg_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  state_reg_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  state_reg_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  state_reg_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  state_reg_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  state_reg_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  state_reg_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  state_reg_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  state_reg_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  state_reg_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  state_reg_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  state_reg_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  state_reg_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  state_reg_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  state_reg_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  state_reg_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  state_pc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  state_csr_misa = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  state_csr_mvendorid = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  state_csr_marchid = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  state_csr_mimpid = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  state_csr_mhartid = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  state_csr_mstatus = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  state_csr_mstatush = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  state_csr_mscratch = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  state_csr_mtvec = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  state_csr_mcounteren = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  state_csr_medeleg = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  state_csr_mideleg = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  state_csr_mip = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  state_csr_mie = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  state_csr_mepc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  state_csr_mcause = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  state_csr_mtval = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  state_csr_cycle = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  state_csr_scounteren = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  state_csr_scause = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  state_csr_stvec = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  state_csr_sepc = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  state_csr_stval = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  state_csr_sscratch = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  state_csr_satp = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  state_csr_pmpcfg0 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  state_csr_pmpcfg1 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  state_csr_pmpcfg2 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  state_csr_pmpcfg3 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  state_csr_pmpaddr0 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  state_csr_pmpaddr1 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  state_csr_pmpaddr2 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  state_csr_pmpaddr3 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  state_csr_MXLEN = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  state_csr_IALIGN = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  state_csr_ILEN = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  state_internal_privilegeMode = _RAND_69[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CheckerWithResult(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mstatush, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_medeleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mideleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_cycle, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_scounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_scause, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_stvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_sepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_stval, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_sscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_satp, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg0, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg1, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg2, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg3, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr0, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr1, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr2, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr3, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [7:0]  io_result_csr_MXLEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [7:0]  io_result_csr_IALIGN, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [7:0]  io_result_csr_ILEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [1:0]  io_result_internal_privilegeMode, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_write_data // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
);
  wire  specCore_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_iFetchpc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [5:0] specCore_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [5:0] specCore_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_now_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [1:0] specCore_io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [1:0] specCore_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  _T = io_mem_read_valid == specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 129:46]
  wire  _T_1 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
  wire  _T_2 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
  wire  _T_3 = ~(io_mem_read_valid == specCore_io_mem_read_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
  wire  _T_4 = io_mem_read_valid | specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 130:43]
  wire  _T_5 = io_mem_read_addr == specCore_io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:47]
  wire  _T_6 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _T_7 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _T_8 = ~(io_mem_read_addr == specCore_io_mem_read_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _T_9 = io_mem_read_memWidth == specCore_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:51]
  wire  _T_10 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _T_11 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _T_12 = ~(io_mem_read_memWidth == specCore_io_mem_read_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _T_13 = io_mem_write_valid == specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 134:47]
  wire  _T_14 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
  wire  _T_15 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
  wire  _T_16 = ~(io_mem_write_valid == specCore_io_mem_write_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
  wire  _T_17 = io_mem_write_valid | specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 135:44]
  wire  _T_18 = io_mem_write_addr == specCore_io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:48]
  wire  _T_19 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _T_20 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _T_21 = ~(io_mem_write_addr == specCore_io_mem_write_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _T_22 = io_mem_write_data == specCore_io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:48]
  wire  _T_23 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _T_24 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _T_25 = ~(io_mem_write_data == specCore_io_mem_write_data); // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _T_26 = io_mem_write_memWidth == specCore_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:52]
  wire  _T_27 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _T_28 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _T_29 = ~(io_mem_write_memWidth == specCore_io_mem_write_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _T_30 = io_instCommit_pc == specCore_io_now_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:39]
  wire  _T_31 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _T_32 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _T_33 = ~(io_instCommit_pc == specCore_io_now_pc); // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _T_34 = io_result_csr_misa == specCore_io_next_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_35 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_36 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_37 = ~(io_result_csr_misa == specCore_io_next_csr_misa); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_38 = io_result_csr_mvendorid == specCore_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_39 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_40 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_41 = ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_42 = io_result_csr_marchid == specCore_io_next_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_43 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_44 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_45 = ~(io_result_csr_marchid == specCore_io_next_csr_marchid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_46 = io_result_csr_mimpid == specCore_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_47 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_48 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_49 = ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_50 = io_result_csr_mhartid == specCore_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_51 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_52 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_53 = ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_54 = io_result_csr_mstatus == specCore_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_55 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_56 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_57 = ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_58 = io_result_csr_mscratch == specCore_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_59 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_60 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_61 = ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_62 = io_result_csr_mtvec == specCore_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_63 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_64 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_65 = ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_66 = io_result_csr_mcounteren == specCore_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_67 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_68 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_69 = ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_70 = io_result_csr_mip == specCore_io_next_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_71 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_72 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_73 = ~(io_result_csr_mip == specCore_io_next_csr_mip); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_74 = io_result_csr_mie == specCore_io_next_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_75 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_76 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_77 = ~(io_result_csr_mie == specCore_io_next_csr_mie); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_78 = io_result_csr_mepc == specCore_io_next_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_79 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_80 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_81 = ~(io_result_csr_mepc == specCore_io_next_csr_mepc); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_82 = io_result_csr_mcause == specCore_io_next_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_83 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_84 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_85 = ~(io_result_csr_mcause == specCore_io_next_csr_mcause); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_86 = io_result_csr_mtval == specCore_io_next_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_87 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_88 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_89 = ~(io_result_csr_mtval == specCore_io_next_csr_mtval); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_90 = io_result_reg_0 == specCore_io_next_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_91 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_92 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_93 = ~(io_result_reg_0 == specCore_io_next_reg_0); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_94 = io_result_reg_1 == specCore_io_next_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_95 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_96 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_97 = ~(io_result_reg_1 == specCore_io_next_reg_1); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_98 = io_result_reg_2 == specCore_io_next_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_99 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_100 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_101 = ~(io_result_reg_2 == specCore_io_next_reg_2); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_102 = io_result_reg_3 == specCore_io_next_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_103 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_104 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_105 = ~(io_result_reg_3 == specCore_io_next_reg_3); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_106 = io_result_reg_4 == specCore_io_next_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_107 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_108 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_109 = ~(io_result_reg_4 == specCore_io_next_reg_4); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_110 = io_result_reg_5 == specCore_io_next_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_111 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_112 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_113 = ~(io_result_reg_5 == specCore_io_next_reg_5); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_114 = io_result_reg_6 == specCore_io_next_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_115 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_116 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_117 = ~(io_result_reg_6 == specCore_io_next_reg_6); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_118 = io_result_reg_7 == specCore_io_next_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_119 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_120 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_121 = ~(io_result_reg_7 == specCore_io_next_reg_7); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_122 = io_result_reg_8 == specCore_io_next_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_123 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_124 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_125 = ~(io_result_reg_8 == specCore_io_next_reg_8); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_126 = io_result_reg_9 == specCore_io_next_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_127 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_128 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_129 = ~(io_result_reg_9 == specCore_io_next_reg_9); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_130 = io_result_reg_10 == specCore_io_next_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_131 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_132 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_133 = ~(io_result_reg_10 == specCore_io_next_reg_10); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_134 = io_result_reg_11 == specCore_io_next_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_135 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_136 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_137 = ~(io_result_reg_11 == specCore_io_next_reg_11); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_138 = io_result_reg_12 == specCore_io_next_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_139 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_140 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_141 = ~(io_result_reg_12 == specCore_io_next_reg_12); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_142 = io_result_reg_13 == specCore_io_next_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_143 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_144 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_145 = ~(io_result_reg_13 == specCore_io_next_reg_13); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_146 = io_result_reg_14 == specCore_io_next_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_147 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_148 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_149 = ~(io_result_reg_14 == specCore_io_next_reg_14); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_150 = io_result_reg_15 == specCore_io_next_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_151 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_152 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_153 = ~(io_result_reg_15 == specCore_io_next_reg_15); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_154 = io_result_reg_16 == specCore_io_next_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_155 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_156 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_157 = ~(io_result_reg_16 == specCore_io_next_reg_16); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_158 = io_result_reg_17 == specCore_io_next_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_159 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_160 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_161 = ~(io_result_reg_17 == specCore_io_next_reg_17); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_162 = io_result_reg_18 == specCore_io_next_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_163 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_164 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_165 = ~(io_result_reg_18 == specCore_io_next_reg_18); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_166 = io_result_reg_19 == specCore_io_next_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_167 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_168 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_169 = ~(io_result_reg_19 == specCore_io_next_reg_19); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_170 = io_result_reg_20 == specCore_io_next_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_171 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_172 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_173 = ~(io_result_reg_20 == specCore_io_next_reg_20); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_174 = io_result_reg_21 == specCore_io_next_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_175 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_176 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_177 = ~(io_result_reg_21 == specCore_io_next_reg_21); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_178 = io_result_reg_22 == specCore_io_next_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_179 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_180 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_181 = ~(io_result_reg_22 == specCore_io_next_reg_22); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_182 = io_result_reg_23 == specCore_io_next_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_183 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_184 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_185 = ~(io_result_reg_23 == specCore_io_next_reg_23); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_186 = io_result_reg_24 == specCore_io_next_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_187 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_188 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_189 = ~(io_result_reg_24 == specCore_io_next_reg_24); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_190 = io_result_reg_25 == specCore_io_next_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_191 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_192 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_193 = ~(io_result_reg_25 == specCore_io_next_reg_25); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_194 = io_result_reg_26 == specCore_io_next_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_195 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_196 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_197 = ~(io_result_reg_26 == specCore_io_next_reg_26); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_198 = io_result_reg_27 == specCore_io_next_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_199 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_200 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_201 = ~(io_result_reg_27 == specCore_io_next_reg_27); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_202 = io_result_reg_28 == specCore_io_next_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_203 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_204 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_205 = ~(io_result_reg_28 == specCore_io_next_reg_28); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_206 = io_result_reg_29 == specCore_io_next_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_207 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_208 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_209 = ~(io_result_reg_29 == specCore_io_next_reg_29); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_210 = io_result_reg_30 == specCore_io_next_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_211 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_212 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_213 = ~(io_result_reg_30 == specCore_io_next_reg_30); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_214 = io_result_reg_31 == specCore_io_next_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_215 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_216 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_217 = ~(io_result_reg_31 == specCore_io_next_reg_31); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_218 = io_event_valid | specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 239:33]
  wire  _T_219 = io_event_valid == specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 241:32]
  wire  _T_220 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _T_221 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _T_222 = ~_T_219; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _T_223 = io_event_intrNO == 32'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:38]
  wire  _T_224 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _T_225 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _T_226 = ~(io_event_intrNO == 32'h0); // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _T_227 = io_event_cause == specCore_io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:37]
  wire  _T_228 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _T_229 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _T_230 = ~(io_event_cause == specCore_io_event_cause); // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _T_231 = io_event_exceptionPC == specCore_io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:43]
  wire  _T_232 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _T_233 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _T_234 = ~(io_event_exceptionPC == specCore_io_event_exceptionPC); // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _T_235 = io_event_exceptionInst == specCore_io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:45]
  wire  _T_236 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  wire  _T_237 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  wire  _T_238 = ~(io_event_exceptionInst == specCore_io_event_exceptionInst); // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  wire  _GEN_0 = _T_4 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _GEN_1 = _T_4 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _GEN_2 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _GEN_3 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _GEN_4 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _GEN_5 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _GEN_6 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_7 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_8 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_9 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_10 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_11 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_12 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_13 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_14 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_15 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_16 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_17 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_18 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_19 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_20 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_21 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_22 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_23 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_24 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_25 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_26 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_27 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_28 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_29 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_30 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_31 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_32 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_33 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_34 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_35 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_36 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_37 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_38 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_39 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_40 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_41 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_42 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_43 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_44 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_45 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_46 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_47 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_48 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_49 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_50 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_51 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_52 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _GEN_53 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _GEN_54 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _GEN_55 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _GEN_56 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  RiscvCore specCore ( // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
    .clock(specCore_clock),
    .reset(specCore_reset),
    .io_inst(specCore_io_inst),
    .io_valid(specCore_io_valid),
    .io_iFetchpc(specCore_io_iFetchpc),
    .io_mem_read_valid(specCore_io_mem_read_valid),
    .io_mem_read_addr(specCore_io_mem_read_addr),
    .io_mem_read_memWidth(specCore_io_mem_read_memWidth),
    .io_mem_read_data(specCore_io_mem_read_data),
    .io_mem_write_valid(specCore_io_mem_write_valid),
    .io_mem_write_addr(specCore_io_mem_write_addr),
    .io_mem_write_memWidth(specCore_io_mem_write_memWidth),
    .io_mem_write_data(specCore_io_mem_write_data),
    .io_now_reg_0(specCore_io_now_reg_0),
    .io_now_reg_1(specCore_io_now_reg_1),
    .io_now_reg_2(specCore_io_now_reg_2),
    .io_now_reg_3(specCore_io_now_reg_3),
    .io_now_reg_4(specCore_io_now_reg_4),
    .io_now_reg_5(specCore_io_now_reg_5),
    .io_now_reg_6(specCore_io_now_reg_6),
    .io_now_reg_7(specCore_io_now_reg_7),
    .io_now_reg_8(specCore_io_now_reg_8),
    .io_now_reg_9(specCore_io_now_reg_9),
    .io_now_reg_10(specCore_io_now_reg_10),
    .io_now_reg_11(specCore_io_now_reg_11),
    .io_now_reg_12(specCore_io_now_reg_12),
    .io_now_reg_13(specCore_io_now_reg_13),
    .io_now_reg_14(specCore_io_now_reg_14),
    .io_now_reg_15(specCore_io_now_reg_15),
    .io_now_reg_16(specCore_io_now_reg_16),
    .io_now_reg_17(specCore_io_now_reg_17),
    .io_now_reg_18(specCore_io_now_reg_18),
    .io_now_reg_19(specCore_io_now_reg_19),
    .io_now_reg_20(specCore_io_now_reg_20),
    .io_now_reg_21(specCore_io_now_reg_21),
    .io_now_reg_22(specCore_io_now_reg_22),
    .io_now_reg_23(specCore_io_now_reg_23),
    .io_now_reg_24(specCore_io_now_reg_24),
    .io_now_reg_25(specCore_io_now_reg_25),
    .io_now_reg_26(specCore_io_now_reg_26),
    .io_now_reg_27(specCore_io_now_reg_27),
    .io_now_reg_28(specCore_io_now_reg_28),
    .io_now_reg_29(specCore_io_now_reg_29),
    .io_now_reg_30(specCore_io_now_reg_30),
    .io_now_reg_31(specCore_io_now_reg_31),
    .io_now_pc(specCore_io_now_pc),
    .io_now_csr_misa(specCore_io_now_csr_misa),
    .io_now_csr_mvendorid(specCore_io_now_csr_mvendorid),
    .io_now_csr_marchid(specCore_io_now_csr_marchid),
    .io_now_csr_mimpid(specCore_io_now_csr_mimpid),
    .io_now_csr_mhartid(specCore_io_now_csr_mhartid),
    .io_now_csr_mstatus(specCore_io_now_csr_mstatus),
    .io_now_csr_mstatush(specCore_io_now_csr_mstatush),
    .io_now_csr_mscratch(specCore_io_now_csr_mscratch),
    .io_now_csr_mtvec(specCore_io_now_csr_mtvec),
    .io_now_csr_mcounteren(specCore_io_now_csr_mcounteren),
    .io_now_csr_medeleg(specCore_io_now_csr_medeleg),
    .io_now_csr_mideleg(specCore_io_now_csr_mideleg),
    .io_now_csr_mip(specCore_io_now_csr_mip),
    .io_now_csr_mie(specCore_io_now_csr_mie),
    .io_now_csr_mepc(specCore_io_now_csr_mepc),
    .io_now_csr_mcause(specCore_io_now_csr_mcause),
    .io_now_csr_mtval(specCore_io_now_csr_mtval),
    .io_now_csr_cycle(specCore_io_now_csr_cycle),
    .io_now_csr_scounteren(specCore_io_now_csr_scounteren),
    .io_now_csr_scause(specCore_io_now_csr_scause),
    .io_now_csr_stvec(specCore_io_now_csr_stvec),
    .io_now_csr_sepc(specCore_io_now_csr_sepc),
    .io_now_csr_stval(specCore_io_now_csr_stval),
    .io_now_csr_sscratch(specCore_io_now_csr_sscratch),
    .io_now_csr_satp(specCore_io_now_csr_satp),
    .io_now_csr_pmpcfg0(specCore_io_now_csr_pmpcfg0),
    .io_now_csr_pmpcfg1(specCore_io_now_csr_pmpcfg1),
    .io_now_csr_pmpcfg2(specCore_io_now_csr_pmpcfg2),
    .io_now_csr_pmpcfg3(specCore_io_now_csr_pmpcfg3),
    .io_now_csr_pmpaddr0(specCore_io_now_csr_pmpaddr0),
    .io_now_csr_pmpaddr1(specCore_io_now_csr_pmpaddr1),
    .io_now_csr_pmpaddr2(specCore_io_now_csr_pmpaddr2),
    .io_now_csr_pmpaddr3(specCore_io_now_csr_pmpaddr3),
    .io_now_csr_MXLEN(specCore_io_now_csr_MXLEN),
    .io_now_csr_IALIGN(specCore_io_now_csr_IALIGN),
    .io_now_csr_ILEN(specCore_io_now_csr_ILEN),
    .io_now_internal_privilegeMode(specCore_io_now_internal_privilegeMode),
    .io_next_reg_0(specCore_io_next_reg_0),
    .io_next_reg_1(specCore_io_next_reg_1),
    .io_next_reg_2(specCore_io_next_reg_2),
    .io_next_reg_3(specCore_io_next_reg_3),
    .io_next_reg_4(specCore_io_next_reg_4),
    .io_next_reg_5(specCore_io_next_reg_5),
    .io_next_reg_6(specCore_io_next_reg_6),
    .io_next_reg_7(specCore_io_next_reg_7),
    .io_next_reg_8(specCore_io_next_reg_8),
    .io_next_reg_9(specCore_io_next_reg_9),
    .io_next_reg_10(specCore_io_next_reg_10),
    .io_next_reg_11(specCore_io_next_reg_11),
    .io_next_reg_12(specCore_io_next_reg_12),
    .io_next_reg_13(specCore_io_next_reg_13),
    .io_next_reg_14(specCore_io_next_reg_14),
    .io_next_reg_15(specCore_io_next_reg_15),
    .io_next_reg_16(specCore_io_next_reg_16),
    .io_next_reg_17(specCore_io_next_reg_17),
    .io_next_reg_18(specCore_io_next_reg_18),
    .io_next_reg_19(specCore_io_next_reg_19),
    .io_next_reg_20(specCore_io_next_reg_20),
    .io_next_reg_21(specCore_io_next_reg_21),
    .io_next_reg_22(specCore_io_next_reg_22),
    .io_next_reg_23(specCore_io_next_reg_23),
    .io_next_reg_24(specCore_io_next_reg_24),
    .io_next_reg_25(specCore_io_next_reg_25),
    .io_next_reg_26(specCore_io_next_reg_26),
    .io_next_reg_27(specCore_io_next_reg_27),
    .io_next_reg_28(specCore_io_next_reg_28),
    .io_next_reg_29(specCore_io_next_reg_29),
    .io_next_reg_30(specCore_io_next_reg_30),
    .io_next_reg_31(specCore_io_next_reg_31),
    .io_next_pc(specCore_io_next_pc),
    .io_next_csr_misa(specCore_io_next_csr_misa),
    .io_next_csr_mvendorid(specCore_io_next_csr_mvendorid),
    .io_next_csr_marchid(specCore_io_next_csr_marchid),
    .io_next_csr_mimpid(specCore_io_next_csr_mimpid),
    .io_next_csr_mhartid(specCore_io_next_csr_mhartid),
    .io_next_csr_mstatus(specCore_io_next_csr_mstatus),
    .io_next_csr_mstatush(specCore_io_next_csr_mstatush),
    .io_next_csr_mscratch(specCore_io_next_csr_mscratch),
    .io_next_csr_mtvec(specCore_io_next_csr_mtvec),
    .io_next_csr_mcounteren(specCore_io_next_csr_mcounteren),
    .io_next_csr_medeleg(specCore_io_next_csr_medeleg),
    .io_next_csr_mideleg(specCore_io_next_csr_mideleg),
    .io_next_csr_mip(specCore_io_next_csr_mip),
    .io_next_csr_mie(specCore_io_next_csr_mie),
    .io_next_csr_mepc(specCore_io_next_csr_mepc),
    .io_next_csr_mcause(specCore_io_next_csr_mcause),
    .io_next_csr_mtval(specCore_io_next_csr_mtval),
    .io_next_csr_cycle(specCore_io_next_csr_cycle),
    .io_next_csr_scounteren(specCore_io_next_csr_scounteren),
    .io_next_csr_scause(specCore_io_next_csr_scause),
    .io_next_csr_stvec(specCore_io_next_csr_stvec),
    .io_next_csr_sepc(specCore_io_next_csr_sepc),
    .io_next_csr_stval(specCore_io_next_csr_stval),
    .io_next_csr_sscratch(specCore_io_next_csr_sscratch),
    .io_next_csr_satp(specCore_io_next_csr_satp),
    .io_next_csr_pmpcfg0(specCore_io_next_csr_pmpcfg0),
    .io_next_csr_pmpcfg1(specCore_io_next_csr_pmpcfg1),
    .io_next_csr_pmpcfg2(specCore_io_next_csr_pmpcfg2),
    .io_next_csr_pmpcfg3(specCore_io_next_csr_pmpcfg3),
    .io_next_csr_pmpaddr0(specCore_io_next_csr_pmpaddr0),
    .io_next_csr_pmpaddr1(specCore_io_next_csr_pmpaddr1),
    .io_next_csr_pmpaddr2(specCore_io_next_csr_pmpaddr2),
    .io_next_csr_pmpaddr3(specCore_io_next_csr_pmpaddr3),
    .io_next_csr_MXLEN(specCore_io_next_csr_MXLEN),
    .io_next_csr_IALIGN(specCore_io_next_csr_IALIGN),
    .io_next_csr_ILEN(specCore_io_next_csr_ILEN),
    .io_next_internal_privilegeMode(specCore_io_next_internal_privilegeMode),
    .io_event_valid(specCore_io_event_valid),
    .io_event_intrNO(specCore_io_event_intrNO),
    .io_event_cause(specCore_io_event_cause),
    .io_event_exceptionPC(specCore_io_event_exceptionPC),
    .io_event_exceptionInst(specCore_io_event_exceptionInst)
  );
  assign specCore_clock = clock;
  assign specCore_reset = reset;
  assign specCore_io_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 116:21]
  assign specCore_io_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 115:21]
  assign specCore_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 140:33]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_mem_read_valid == specCore_io_mem_read_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:129 assert(regDelay(io.mem.get.read.valid) === regDelay(specCore.io.mem.read.valid))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & _T_2 & ~(io_mem_read_addr == specCore_io_mem_read_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:131 assert(regDelay(io.mem.get.read.addr) === regDelay(specCore.io.mem.read.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_0 & ~(io_mem_read_memWidth == specCore_io_mem_read_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:132 assert(regDelay(io.mem.get.read.memWidth) === regDelay(specCore.io.mem.read.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(io_mem_write_valid == specCore_io_mem_write_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:134 assert(regDelay(io.mem.get.write.valid) === regDelay(specCore.io.mem.write.valid))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17 & _T_2 & ~(io_mem_write_addr == specCore_io_mem_write_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:136 assert(regDelay(io.mem.get.write.addr) === regDelay(specCore.io.mem.write.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2 & ~(io_mem_write_data == specCore_io_mem_write_data)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:137 assert(regDelay(io.mem.get.write.data) === regDelay(specCore.io.mem.write.data))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2 & ~(io_mem_write_memWidth == specCore_io_mem_write_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:138 assert(regDelay(io.mem.get.write.memWidth) === regDelay(specCore.io.mem.write.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_instCommit_valid & _T_2 & ~(io_instCommit_pc == specCore_io_now_pc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:225 assert(regDelay(io.instCommit.pc) === regDelay(specCore.io.now.pc))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_misa == specCore_io_next_csr_misa)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_marchid == specCore_io_next_csr_marchid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mip == specCore_io_next_csr_mip)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mie == specCore_io_next_csr_mie)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mepc == specCore_io_next_csr_mepc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mcause == specCore_io_next_csr_mcause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mtval == specCore_io_next_csr_mtval)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_0 == specCore_io_next_reg_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_1 == specCore_io_next_reg_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_2 == specCore_io_next_reg_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_3 == specCore_io_next_reg_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_4 == specCore_io_next_reg_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_5 == specCore_io_next_reg_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_6 == specCore_io_next_reg_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_7 == specCore_io_next_reg_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_8 == specCore_io_next_reg_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_9 == specCore_io_next_reg_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_10 == specCore_io_next_reg_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_11 == specCore_io_next_reg_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_12 == specCore_io_next_reg_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_13 == specCore_io_next_reg_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_14 == specCore_io_next_reg_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_15 == specCore_io_next_reg_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_16 == specCore_io_next_reg_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_17 == specCore_io_next_reg_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_18 == specCore_io_next_reg_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_19 == specCore_io_next_reg_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_20 == specCore_io_next_reg_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_21 == specCore_io_next_reg_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_22 == specCore_io_next_reg_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_23 == specCore_io_next_reg_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_24 == specCore_io_next_reg_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_25 == specCore_io_next_reg_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_26 == specCore_io_next_reg_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_27 == specCore_io_next_reg_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_28 == specCore_io_next_reg_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_29 == specCore_io_next_reg_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_30 == specCore_io_next_reg_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_31 == specCore_io_next_reg_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_218 & _T_2 & ~_T_219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Checker.scala:240 assert(\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_intrNO == 32'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:243 assert(regDelay(io.event.intrNO) === regDelay(specCore.io.event.intrNO))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_cause == specCore_io_event_cause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:244 assert(regDelay(io.event.cause) === regDelay(specCore.io.event.cause))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_exceptionPC == specCore_io_event_exceptionPC)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:245 assert(regDelay(io.event.exceptionPC) === regDelay(specCore.io.event.exceptionPC))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_exceptionInst == specCore_io_event_exceptionInst)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:246 assert(regDelay(io.event.exceptionInst) === regDelay(specCore.io.event.exceptionInst))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(io_mem_read_valid == specCore_io_mem_read_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_mem_read_addr == specCore_io_mem_read_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_mem_read_memWidth == specCore_io_mem_read_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
    end
    //
    if (_T_2) begin
      assert(io_mem_write_valid == specCore_io_mem_write_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
    end
    //
    if (_T_17 & _T_2) begin
      assert(io_mem_write_addr == specCore_io_mem_write_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
    end
    //
    if (_T_17 & _T_2) begin
      assert(io_mem_write_data == specCore_io_mem_write_data); // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
    end
    //
    if (_T_17 & _T_2) begin
      assert(io_mem_write_memWidth == specCore_io_mem_write_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_instCommit_pc == specCore_io_now_pc); // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_misa == specCore_io_next_csr_misa); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_marchid == specCore_io_next_csr_marchid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mimpid == specCore_io_next_csr_mimpid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mhartid == specCore_io_next_csr_mhartid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mstatus == specCore_io_next_csr_mstatus); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mscratch == specCore_io_next_csr_mscratch); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mtvec == specCore_io_next_csr_mtvec); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mip == specCore_io_next_csr_mip); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mie == specCore_io_next_csr_mie); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mepc == specCore_io_next_csr_mepc); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mcause == specCore_io_next_csr_mcause); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mtval == specCore_io_next_csr_mtval); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_0 == specCore_io_next_reg_0); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_1 == specCore_io_next_reg_1); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_2 == specCore_io_next_reg_2); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_3 == specCore_io_next_reg_3); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_4 == specCore_io_next_reg_4); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_5 == specCore_io_next_reg_5); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_6 == specCore_io_next_reg_6); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_7 == specCore_io_next_reg_7); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_8 == specCore_io_next_reg_8); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_9 == specCore_io_next_reg_9); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_10 == specCore_io_next_reg_10); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_11 == specCore_io_next_reg_11); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_12 == specCore_io_next_reg_12); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_13 == specCore_io_next_reg_13); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_14 == specCore_io_next_reg_14); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_15 == specCore_io_next_reg_15); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_16 == specCore_io_next_reg_16); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_17 == specCore_io_next_reg_17); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_18 == specCore_io_next_reg_18); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_19 == specCore_io_next_reg_19); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_20 == specCore_io_next_reg_20); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_21 == specCore_io_next_reg_21); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_22 == specCore_io_next_reg_22); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_23 == specCore_io_next_reg_23); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_24 == specCore_io_next_reg_24); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_25 == specCore_io_next_reg_25); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_26 == specCore_io_next_reg_26); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_27 == specCore_io_next_reg_27); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_28 == specCore_io_next_reg_28); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_29 == specCore_io_next_reg_29); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_30 == specCore_io_next_reg_30); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_31 == specCore_io_next_reg_31); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (_T_218 & _T_2) begin
      assert(_T_219); // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_intrNO == 32'h0); // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_cause == specCore_io_event_cause); // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_exceptionPC == specCore_io_event_exceptionPC); // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_exceptionInst == specCore_io_event_exceptionInst); // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
    end
  end
endmodule
module CheckerWrapper(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mstatush, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_medeleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mideleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_cycle, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_scounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_scause, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_stvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_sepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_stval, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_sscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_satp, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg0, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg1, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg2, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg3, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr0, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr1, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr2, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr3, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [7:0]  io_result_csr_MXLEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [7:0]  io_result_csr_IALIGN, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [7:0]  io_result_csr_ILEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [1:0]  io_result_internal_privilegeMode, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_write_data // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
);
  wire  checker__clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_instCommit_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [7:0] checker__io_result_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [7:0] checker__io_result_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [7:0] checker__io_result_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [1:0] checker__io_result_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [5:0] checker__io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [5:0] checker__io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  CheckerWithResult checker_ ( // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
    .clock(checker__clock),
    .reset(checker__reset),
    .io_instCommit_valid(checker__io_instCommit_valid),
    .io_instCommit_inst(checker__io_instCommit_inst),
    .io_instCommit_pc(checker__io_instCommit_pc),
    .io_result_reg_0(checker__io_result_reg_0),
    .io_result_reg_1(checker__io_result_reg_1),
    .io_result_reg_2(checker__io_result_reg_2),
    .io_result_reg_3(checker__io_result_reg_3),
    .io_result_reg_4(checker__io_result_reg_4),
    .io_result_reg_5(checker__io_result_reg_5),
    .io_result_reg_6(checker__io_result_reg_6),
    .io_result_reg_7(checker__io_result_reg_7),
    .io_result_reg_8(checker__io_result_reg_8),
    .io_result_reg_9(checker__io_result_reg_9),
    .io_result_reg_10(checker__io_result_reg_10),
    .io_result_reg_11(checker__io_result_reg_11),
    .io_result_reg_12(checker__io_result_reg_12),
    .io_result_reg_13(checker__io_result_reg_13),
    .io_result_reg_14(checker__io_result_reg_14),
    .io_result_reg_15(checker__io_result_reg_15),
    .io_result_reg_16(checker__io_result_reg_16),
    .io_result_reg_17(checker__io_result_reg_17),
    .io_result_reg_18(checker__io_result_reg_18),
    .io_result_reg_19(checker__io_result_reg_19),
    .io_result_reg_20(checker__io_result_reg_20),
    .io_result_reg_21(checker__io_result_reg_21),
    .io_result_reg_22(checker__io_result_reg_22),
    .io_result_reg_23(checker__io_result_reg_23),
    .io_result_reg_24(checker__io_result_reg_24),
    .io_result_reg_25(checker__io_result_reg_25),
    .io_result_reg_26(checker__io_result_reg_26),
    .io_result_reg_27(checker__io_result_reg_27),
    .io_result_reg_28(checker__io_result_reg_28),
    .io_result_reg_29(checker__io_result_reg_29),
    .io_result_reg_30(checker__io_result_reg_30),
    .io_result_reg_31(checker__io_result_reg_31),
    .io_result_pc(checker__io_result_pc),
    .io_result_csr_misa(checker__io_result_csr_misa),
    .io_result_csr_mvendorid(checker__io_result_csr_mvendorid),
    .io_result_csr_marchid(checker__io_result_csr_marchid),
    .io_result_csr_mimpid(checker__io_result_csr_mimpid),
    .io_result_csr_mhartid(checker__io_result_csr_mhartid),
    .io_result_csr_mstatus(checker__io_result_csr_mstatus),
    .io_result_csr_mstatush(checker__io_result_csr_mstatush),
    .io_result_csr_mscratch(checker__io_result_csr_mscratch),
    .io_result_csr_mtvec(checker__io_result_csr_mtvec),
    .io_result_csr_mcounteren(checker__io_result_csr_mcounteren),
    .io_result_csr_medeleg(checker__io_result_csr_medeleg),
    .io_result_csr_mideleg(checker__io_result_csr_mideleg),
    .io_result_csr_mip(checker__io_result_csr_mip),
    .io_result_csr_mie(checker__io_result_csr_mie),
    .io_result_csr_mepc(checker__io_result_csr_mepc),
    .io_result_csr_mcause(checker__io_result_csr_mcause),
    .io_result_csr_mtval(checker__io_result_csr_mtval),
    .io_result_csr_cycle(checker__io_result_csr_cycle),
    .io_result_csr_scounteren(checker__io_result_csr_scounteren),
    .io_result_csr_scause(checker__io_result_csr_scause),
    .io_result_csr_stvec(checker__io_result_csr_stvec),
    .io_result_csr_sepc(checker__io_result_csr_sepc),
    .io_result_csr_stval(checker__io_result_csr_stval),
    .io_result_csr_sscratch(checker__io_result_csr_sscratch),
    .io_result_csr_satp(checker__io_result_csr_satp),
    .io_result_csr_pmpcfg0(checker__io_result_csr_pmpcfg0),
    .io_result_csr_pmpcfg1(checker__io_result_csr_pmpcfg1),
    .io_result_csr_pmpcfg2(checker__io_result_csr_pmpcfg2),
    .io_result_csr_pmpcfg3(checker__io_result_csr_pmpcfg3),
    .io_result_csr_pmpaddr0(checker__io_result_csr_pmpaddr0),
    .io_result_csr_pmpaddr1(checker__io_result_csr_pmpaddr1),
    .io_result_csr_pmpaddr2(checker__io_result_csr_pmpaddr2),
    .io_result_csr_pmpaddr3(checker__io_result_csr_pmpaddr3),
    .io_result_csr_MXLEN(checker__io_result_csr_MXLEN),
    .io_result_csr_IALIGN(checker__io_result_csr_IALIGN),
    .io_result_csr_ILEN(checker__io_result_csr_ILEN),
    .io_result_internal_privilegeMode(checker__io_result_internal_privilegeMode),
    .io_event_valid(checker__io_event_valid),
    .io_event_intrNO(checker__io_event_intrNO),
    .io_event_cause(checker__io_event_cause),
    .io_event_exceptionPC(checker__io_event_exceptionPC),
    .io_event_exceptionInst(checker__io_event_exceptionInst),
    .io_mem_read_valid(checker__io_mem_read_valid),
    .io_mem_read_addr(checker__io_mem_read_addr),
    .io_mem_read_memWidth(checker__io_mem_read_memWidth),
    .io_mem_read_data(checker__io_mem_read_data),
    .io_mem_write_valid(checker__io_mem_write_valid),
    .io_mem_write_addr(checker__io_mem_write_addr),
    .io_mem_write_memWidth(checker__io_mem_write_memWidth),
    .io_mem_write_data(checker__io_mem_write_data)
  );
  assign checker__clock = clock;
  assign checker__reset = reset;
  assign checker__io_instCommit_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 361:25]
  assign checker__io_instCommit_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 361:25]
  assign checker__io_instCommit_pc = io_instCommit_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 361:25]
  assign checker__io_result_reg_0 = io_result_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_1 = io_result_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_2 = io_result_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_3 = io_result_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_4 = io_result_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_5 = io_result_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_6 = io_result_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_7 = io_result_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_8 = io_result_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_9 = io_result_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_10 = io_result_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_11 = io_result_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_12 = io_result_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_13 = io_result_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_14 = io_result_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_15 = io_result_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_16 = io_result_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_17 = io_result_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_18 = io_result_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_19 = io_result_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_20 = io_result_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_21 = io_result_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_22 = io_result_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_23 = io_result_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_24 = io_result_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_25 = io_result_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_26 = io_result_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_27 = io_result_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_28 = io_result_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_29 = io_result_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_30 = io_result_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_31 = io_result_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_pc = io_result_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_misa = io_result_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mvendorid = io_result_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_marchid = io_result_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mimpid = io_result_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mhartid = io_result_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mstatus = io_result_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mstatush = io_result_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mscratch = io_result_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mtvec = io_result_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mcounteren = io_result_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_medeleg = io_result_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mideleg = io_result_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mip = io_result_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mie = io_result_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mepc = io_result_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mcause = io_result_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mtval = io_result_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_cycle = io_result_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_scounteren = io_result_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_scause = io_result_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_stvec = io_result_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_sepc = io_result_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_stval = io_result_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_sscratch = io_result_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_satp = io_result_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg0 = io_result_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg1 = io_result_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg2 = io_result_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg3 = io_result_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr0 = io_result_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr1 = io_result_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr2 = io_result_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr3 = io_result_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_MXLEN = io_result_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_IALIGN = io_result_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_ILEN = io_result_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_internal_privilegeMode = io_result_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_event_valid = io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_intrNO = io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_cause = io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_exceptionPC = io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_exceptionInst = io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_mem_read_valid = io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_read_addr = io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_read_memWidth = io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_valid = io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_addr = io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_memWidth = io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_data = io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
endmodule
