`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  wire [0:0] PI_clock = clock;
  reg [0:0] PI_reset;
  top_formal UUT (
    .clock(PI_clock),
    .reset(PI_reset)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$11525  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$11555  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$11837  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$11855  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:101:execute$11861  = 1'b0;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11529  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11535  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11541  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11547  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11553  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11559  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11565  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11571  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11577  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11583  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11589  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11595  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11601  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11607  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11613  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11619  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11625  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11631  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11637  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11643  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11649  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11655  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11661  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11667  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11673  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11679  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11685  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11691  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11697  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11703  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11709  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11715  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11721  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11727  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11733  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11739  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11745  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11751  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11757  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11763  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11769  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11775  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11781  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11787  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11793  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11799  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11805  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11811  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11817  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11823  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11829  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11835  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11841  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11847  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11853  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11859  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11865  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11871  = 1'b1;
    // UUT.checker_inst.checker_.$auto$async2sync.\cc:110:execute$11877  = 1'b1;
    UUT.checker_inst.checker_.specCore.state_csr_IALIGN = 8'b00000000;
    UUT.checker_inst.checker_.specCore.state_csr_ILEN = 8'b00000000;
    UUT.checker_inst.checker_.specCore.state_csr_MXLEN = 8'b00000000;
    UUT.checker_inst.checker_.specCore.state_csr_cycle = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_marchid = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mcause = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mcounteren = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_medeleg = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mepc = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mhartid = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mideleg = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mie = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mimpid = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mip = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_misa = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mscratch = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mstatus = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mstatush = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mtval = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mtvec = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_mvendorid = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpaddr0 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpaddr1 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpaddr2 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpaddr3 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpcfg0 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpcfg1 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpcfg2 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_pmpcfg3 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_satp = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_scause = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_scounteren = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_sepc = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_sscratch = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_stval = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_csr_stvec = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_internal_privilegeMode = 2'b00;
    UUT.checker_inst.checker_.specCore.state_pc = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_0 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_1 = 32'b01111111111111111111111111111100;
    UUT.checker_inst.checker_.specCore.state_reg_10 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_11 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_12 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_13 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_14 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_15 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_16 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_17 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_18 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_19 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_2 = 32'b01111111111111111111111111111100;
    UUT.checker_inst.checker_.specCore.state_reg_20 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_21 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_22 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_23 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_24 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_25 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_26 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_27 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_28 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_29 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_3 = 32'b00000000000000000111111111111000;
    UUT.checker_inst.checker_.specCore.state_reg_30 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_31 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_4 = 32'b00000000000000010000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_5 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_6 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_7 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_8 = 32'b00000000000000000000000000000000;
    UUT.checker_inst.checker_.specCore.state_reg_9 = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.captured_rmask = 4'b0000;
    UUT.wrapper_inst.captured_wstrb = 4'b0000;
    UUT.wrapper_inst.csr_mcause = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.mem_addr_reg = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.mem_data_reg = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.mem_read_valid_reg = 1'b0;
    UUT.wrapper_inst.mem_write_valid_reg = 1'b0;
    UUT.wrapper_inst.result_csr_mie = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.result_csr_mip = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.result_csr_mstatus = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.result_csr_mstatush = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[10]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[11]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[12]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[13]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[14]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[15]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[16]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[17]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[18]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[19]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[20]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[21]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[22]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[23]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[24]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[25]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[26]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[27]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[28]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[29]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[30]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[31]  = 32'b10000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[4]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[5]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[6]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[7]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[8]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.\shadow_regfile[9]  = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_custom_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_hpm_counter_value = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_hpm_counterh_value = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_hpm_event_value = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mcause_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mepc_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mie_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mip_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_misa_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mscratch_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mstatus_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mstatush_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mtval_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.csr_mtvec_value = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.mem_rd_enable_q = 1'b0;
    UUT.wrapper_inst.uut.mem_rd_func_q = 5'b00000;
    UUT.wrapper_inst.uut.mem_rd_reg_q = 5'b00000;
    UUT.wrapper_inst.uut.mem_wr_enable_q = 1'b0;
    UUT.wrapper_inst.uut.next_rvfi_intr = 1'b0;
    UUT.wrapper_inst.uut.pc = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.reset_q = 1'b0;
    UUT.wrapper_inst.uut.rvfi_csr_custom_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_ro_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_ro_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_ro_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_ro_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_custom_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_marchid_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_marchid_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_marchid_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_marchid_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcause_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcause_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcause_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcause_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mconfigptr_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mconfigptr_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mconfigptr_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mconfigptr_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycle_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycle_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycle_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycle_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycleh_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycleh_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycleh_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mcycleh_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mepc_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mepc_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mepc_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mepc_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhartid_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhartid_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhartid_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhartid_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter10h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter11h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter12h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter13h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter14h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter15h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter16h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter17h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter18h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter19h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter20h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter21h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter22h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter23h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter24h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter25h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter26h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter27h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter28h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter29h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter30h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter31h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter3h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter4h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter5h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter6h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter7h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter8h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9h_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9h_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9h_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmcounter9h_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent10_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent10_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent10_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent10_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent11_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent11_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent11_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent11_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent12_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent12_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent12_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent12_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent13_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent13_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent13_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent13_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent14_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent14_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent14_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent14_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent15_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent15_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent15_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent15_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent16_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent16_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent16_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent16_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent17_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent17_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent17_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent17_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent18_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent18_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent18_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent18_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent19_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent19_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent19_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent19_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent20_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent20_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent20_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent20_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent21_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent21_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent21_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent21_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent22_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent22_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent22_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent22_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent23_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent23_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent23_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent23_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent24_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent24_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent24_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent24_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent25_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent25_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent25_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent25_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent26_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent26_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent26_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent26_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent27_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent27_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent27_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent27_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent28_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent28_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent28_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent28_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent29_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent29_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent29_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent29_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent30_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent30_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent30_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent30_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent31_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent31_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent31_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent31_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent3_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent3_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent3_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent3_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent4_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent4_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent4_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent4_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent5_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent5_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent5_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent5_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent6_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent6_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent6_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent6_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent7_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent7_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent7_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent7_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent8_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent8_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent8_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent8_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent9_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent9_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent9_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mhpmevent9_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mie_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mie_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mie_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mie_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mimpid_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mimpid_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mimpid_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mimpid_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstret_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstret_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstret_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstret_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstreth_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstreth_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstreth_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_minstreth_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mip_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mip_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mip_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mip_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_misa_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_misa_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_misa_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_misa_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mscratch_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mscratch_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mscratch_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mscratch_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatus_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatus_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatus_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatus_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatush_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatush_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatush_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mstatush_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtval_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtval_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtval_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtval_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtvec_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtvec_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtvec_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mtvec_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mvendorid_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mvendorid_rmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mvendorid_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_csr_mvendorid_wmask = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_halt = 1'b0;
    UUT.wrapper_inst.uut.rvfi_insn = 32'b00000000010000000000000000110011;
    UUT.wrapper_inst.uut.rvfi_intr = 1'b0;
    UUT.wrapper_inst.uut.rvfi_ixl = 2'b00;
    UUT.wrapper_inst.uut.rvfi_mem_addr = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_mem_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_mem_rmask = 4'b0000;
    UUT.wrapper_inst.uut.rvfi_mem_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_mem_wmask = 4'b0000;
    UUT.wrapper_inst.uut.rvfi_mode = 2'b00;
    UUT.wrapper_inst.uut.rvfi_order = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_pc_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_pc_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_rd_addr = 5'b00000;
    UUT.wrapper_inst.uut.rvfi_rd_wdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_rs1_addr = 5'b00000;
    UUT.wrapper_inst.uut.rvfi_rs1_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_rs2_addr = 5'b00000;
    UUT.wrapper_inst.uut.rvfi_rs2_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.uut.rvfi_trap = 1'b0;
    UUT.wrapper_inst.uut.rvfi_valid = 1'b1;
    UUT.wrapper_inst.uut.regfile[5'b00000] = 32'b00000000000000000000000000000000;

    // state 0
    PI_reset = 1'b1;
    UUT.wrapper_inst.irq = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.dmem_rdata = 32'b00000000000000000000000000000000;
    UUT.wrapper_inst.stall = 1'b0;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_reset <= 1'b0;
      UUT.wrapper_inst.irq <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.dmem_rdata <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.stall <= 1'b0;
    end

    // state 2
    if (cycle == 1) begin
      PI_reset <= 1'b0;
      UUT.wrapper_inst.irq <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.dmem_rdata <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.stall <= 1'b0;
    end

    // state 3
    if (cycle == 2) begin
      PI_reset <= 1'b0;
      UUT.wrapper_inst.irq <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.dmem_rdata <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.stall <= 1'b0;
    end

    // state 4
    if (cycle == 3) begin
      PI_reset <= 1'b0;
      UUT.wrapper_inst.irq <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.dmem_rdata <= 32'b00000000000000000000000000000000;
      UUT.wrapper_inst.stall <= 1'b0;
    end

    genclock <= cycle < 4;
    cycle <= cycle + 1;
  end
endmodule
