`define SYNTHESIS 
`define NERV_RVFI
`define NERV_CSR