module RiscvTrans(
  input         clock,
  input         reset,
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_iFetchpc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [31:0] io_now_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [1:0]  io_now_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_next_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [1:0]  io_next_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [31:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
);
  wire  _exceptionVec_WIRE_5 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_5 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_7 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_7 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_1 = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_13 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_13 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_2 = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_15 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_15 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_3 = 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] inst = io_valid ? io_inst : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_3257 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _T_426 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_427 = 32'h5003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_444 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _T_614 = inst & 32'hfe007fff; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_615 = 32'h12000073 == _T_614; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_616 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_48 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_608 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_609 = 32'h10500073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_610 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_47 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_601 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_602 = 32'h30200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_603 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_46 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_594 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_595 = 32'h10200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_596 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_45 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_587 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_588 = 32'h2007033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_589 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_590 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_44 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_580 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_581 = 32'h2006033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_582 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_583 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_43 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_573 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_574 = 32'h2005033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_575 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_576 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_42 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_566 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_567 = 32'h2004033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_568 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_569 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_41 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_559 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_560 = 32'h2003033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_561 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_562 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_40 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_552 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_553 = 32'h2002033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_554 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_555 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_39 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_545 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_546 = 32'h2001033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_547 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_548 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_38 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_538 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_539 = 32'h2000033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_540 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_541 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_37 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_532 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_533 = 32'hf == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_534 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_36 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_523 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_524 = 32'h73 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_525 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_35 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_517 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire  _T_518 = 32'h100073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_519 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_34 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_493 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_494 = 32'h2023 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_495 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_496 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_33 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_469 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_470 = 32'h1023 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_471 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_472 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_32 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_446 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_447 = 32'h23 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_448 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_449 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_31 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [19:0] _T_428 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_30 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_407 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_408 = 32'h4003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_409 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_29 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_387 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_388 = 32'h2003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_389 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_28 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_367 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_368 = 32'h1003 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_369 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_27 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_347 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_348 = 32'h3 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_349 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_26 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_320 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_321 = 32'h7063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_322 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_323 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_324 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_25 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_291 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_292 = 32'h5063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_293 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_294 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_295 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_24 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_264 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_265 = 32'h6063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_266 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_267 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_268 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_23 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_235 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_236 = 32'h4063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_237 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_238 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_239 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_22 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_208 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_209 = 32'h1063 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_210 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_211 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_212 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_21 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_181 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_182 = 32'h63 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_183 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [24:0] _T_184 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_185 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_20 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_156 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_157 = 32'h67 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_158 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_19 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_125 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_126 = 32'h40005033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_127 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_128 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_18 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_118 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_119 = 32'h40000033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_120 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_121 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_17 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_111 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_112 = 32'h5033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_113 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_114 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_16 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_104 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_105 = 32'h1033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_106 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_107 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_15 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_97 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_98 = 32'h4033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_99 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_100 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_14 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_90 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_91 = 32'h6033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_92 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_93 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_13 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_83 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_84 = 32'h7033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_85 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_86 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_12 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_76 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_77 = 32'h3033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_78 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_79 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_11 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_69 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_70 = 32'h2033 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_71 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_72 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_10 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_62 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_63 = 32'h33 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [24:0] _T_64 = inst[24:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [19:0] _T_65 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_9 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_48 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_49 = 32'h40005013 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [19:0] _T_50 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_8 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_42 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_43 = 32'h5013 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [19:0] _T_44 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_7 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_36 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_37 = 32'h1013 == _T_587; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [19:0] _T_38 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_6 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_30 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_31 = 32'h4013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_32 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_5 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_24 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_25 = 32'h6013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_26 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_4 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_18 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_19 = 32'h7013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_20 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_3 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_12 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_13 = 32'h3013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_14 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_2 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_6 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_7 = 32'h2013 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_8 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T_1 = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1 = 32'h13 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _T_2 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rs1_T = inst[19:15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_66 = _T_1 ? inst[19:15] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [4:0] _GEN_137 = _T_7 ? inst[19:15] : _GEN_66; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_208 = _T_13 ? inst[19:15] : _GEN_137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_279 = _T_19 ? inst[19:15] : _GEN_208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_350 = _T_25 ? inst[19:15] : _GEN_279; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_421 = _T_31 ? inst[19:15] : _GEN_350; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_492 = _T_37 ? inst[19:15] : _GEN_421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_563 = _T_43 ? inst[19:15] : _GEN_492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_634 = _T_49 ? inst[19:15] : _GEN_563; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_876 = _T_63 ? inst[19:15] : _GEN_634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_947 = _T_70 ? inst[19:15] : _GEN_876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1018 = _T_77 ? inst[19:15] : _GEN_947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1089 = _T_84 ? inst[19:15] : _GEN_1018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1160 = _T_91 ? inst[19:15] : _GEN_1089; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1231 = _T_98 ? inst[19:15] : _GEN_1160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1302 = _T_105 ? inst[19:15] : _GEN_1231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1373 = _T_112 ? inst[19:15] : _GEN_1302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1444 = _T_119 ? inst[19:15] : _GEN_1373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1515 = _T_126 ? inst[19:15] : _GEN_1444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1736 = _T_157 ? inst[19:15] : _GEN_1515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1792 = _T_182 ? inst[19:15] : _GEN_1736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1817 = _T_209 ? inst[19:15] : _GEN_1792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1842 = _T_236 ? inst[19:15] : _GEN_1817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1867 = _T_265 ? inst[19:15] : _GEN_1842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1892 = _T_292 ? inst[19:15] : _GEN_1867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1917 = _T_321 ? inst[19:15] : _GEN_1892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1999 = _T_348 ? inst[19:15] : _GEN_1917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2112 = _T_368 ? inst[19:15] : _GEN_1999; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2225 = _T_388 ? inst[19:15] : _GEN_2112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2303 = _T_408 ? inst[19:15] : _GEN_2225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2416 = _T_427 ? inst[19:15] : _GEN_2303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2463 = _T_447 ? inst[19:15] : _GEN_2416; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2483 = _T_470 ? inst[19:15] : _GEN_2463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2503 = _T_494 ? inst[19:15] : _GEN_2483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2516 = _T_518 ? inst[19:15] : _GEN_2503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2534 = _T_524 ? inst[19:15] : _GEN_2516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2545 = _T_533 ? inst[19:15] : _GEN_2534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2585 = _T_539 ? inst[19:15] : _GEN_2545; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2656 = _T_546 ? inst[19:15] : _GEN_2585; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2727 = _T_553 ? inst[19:15] : _GEN_2656; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2798 = _T_560 ? inst[19:15] : _GEN_2727; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2869 = _T_567 ? inst[19:15] : _GEN_2798; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2940 = _T_574 ? inst[19:15] : _GEN_2869; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3011 = _T_581 ? inst[19:15] : _GEN_2940; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3082 = _T_588 ? inst[19:15] : _GEN_3011; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3131 = _T_595 ? inst[19:15] : _GEN_3082; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3152 = _T_602 ? inst[19:15] : _GEN_3131; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3166 = _T_609 ? inst[19:15] : _GEN_3152; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3173 = _T_615 ? inst[19:15] : _GEN_3166; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs1 = io_valid ? _GEN_3173 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [4:0] _GEN_3260 = rs1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [31:0] now_reg_31 = io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_30 = io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_29 = io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_28 = io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_27 = io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_26 = io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_25 = io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_24 = io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_23 = io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_22 = io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_21 = io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_20 = io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_19 = io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_18 = io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_17 = io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_16 = io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_15 = io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_14 = io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_13 = io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_12 = io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_11 = io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_10 = io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_9 = io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_8 = io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_7 = io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_6 = io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_5 = io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_4 = io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_3 = io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_2 = io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_1 = io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_reg_0 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_0 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_1 = 5'h1 == rs1 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_2 = 5'h2 == rs1 ? io_now_reg_2 : _GEN_1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_3 = 5'h3 == rs1 ? io_now_reg_3 : _GEN_2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_4 = 5'h4 == rs1 ? io_now_reg_4 : _GEN_3; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_5 = 5'h5 == rs1 ? io_now_reg_5 : _GEN_4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_6 = 5'h6 == rs1 ? io_now_reg_6 : _GEN_5; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_7 = 5'h7 == rs1 ? io_now_reg_7 : _GEN_6; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_8 = 5'h8 == rs1 ? io_now_reg_8 : _GEN_7; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_9 = 5'h9 == rs1 ? io_now_reg_9 : _GEN_8; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_10 = 5'ha == rs1 ? io_now_reg_10 : _GEN_9; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_11 = 5'hb == rs1 ? io_now_reg_11 : _GEN_10; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_12 = 5'hc == rs1 ? io_now_reg_12 : _GEN_11; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_13 = 5'hd == rs1 ? io_now_reg_13 : _GEN_12; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_14 = 5'he == rs1 ? io_now_reg_14 : _GEN_13; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_15 = 5'hf == rs1 ? io_now_reg_15 : _GEN_14; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_16 = 5'h10 == rs1 ? io_now_reg_16 : _GEN_15; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_17 = 5'h11 == rs1 ? io_now_reg_17 : _GEN_16; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_18 = 5'h12 == rs1 ? io_now_reg_18 : _GEN_17; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_19 = 5'h13 == rs1 ? io_now_reg_19 : _GEN_18; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_20 = 5'h14 == rs1 ? io_now_reg_20 : _GEN_19; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_21 = 5'h15 == rs1 ? io_now_reg_21 : _GEN_20; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_22 = 5'h16 == rs1 ? io_now_reg_22 : _GEN_21; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_23 = 5'h17 == rs1 ? io_now_reg_23 : _GEN_22; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_24 = 5'h18 == rs1 ? io_now_reg_24 : _GEN_23; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_25 = 5'h19 == rs1 ? io_now_reg_25 : _GEN_24; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_26 = 5'h1a == rs1 ? io_now_reg_26 : _GEN_25; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_27 = 5'h1b == rs1 ? io_now_reg_27 : _GEN_26; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_28 = 5'h1c == rs1 ? io_now_reg_28 : _GEN_27; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_29 = 5'h1d == rs1 ? io_now_reg_29 : _GEN_28; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_30 = 5'h1e == rs1 ? io_now_reg_30 : _GEN_29; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_31 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs1_37 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [11:0] _imm_11_0_T_21 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_20 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_19 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_18 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_17 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_16 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_15 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_14 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_13 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_12 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_11 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_10 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_9 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_8 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_7 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_6 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_5 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_4 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_3 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_2 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T_1 = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _imm_11_0_T = inst[31:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _GEN_65 = _T_1 ? inst[31:20] : 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire [11:0] _GEN_136 = _T_7 ? inst[31:20] : _GEN_65; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_207 = _T_13 ? inst[31:20] : _GEN_136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_278 = _T_19 ? inst[31:20] : _GEN_207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_349 = _T_25 ? inst[31:20] : _GEN_278; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_420 = _T_31 ? inst[31:20] : _GEN_349; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_491 = _T_37 ? inst[31:20] : _GEN_420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_562 = _T_43 ? inst[31:20] : _GEN_491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_633 = _T_49 ? inst[31:20] : _GEN_562; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1735 = _T_157 ? inst[31:20] : _GEN_633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1998 = _T_348 ? inst[31:20] : _GEN_1735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2111 = _T_368 ? inst[31:20] : _GEN_1998; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2224 = _T_388 ? inst[31:20] : _GEN_2111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2302 = _T_408 ? inst[31:20] : _GEN_2224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2415 = _T_427 ? inst[31:20] : _GEN_2302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2515 = _T_518 ? inst[31:20] : _GEN_2415; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2533 = _T_524 ? inst[31:20] : _GEN_2515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2544 = _T_533 ? inst[31:20] : _GEN_2533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3130 = _T_595 ? inst[31:20] : _GEN_2544; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3151 = _T_602 ? inst[31:20] : _GEN_3130; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3165 = _T_609 ? inst[31:20] : _GEN_3151; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3172 = _T_615 ? inst[31:20] : _GEN_3165; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] imm_11_0 = io_valid ? _GEN_3172 : 12'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire [11:0] _GEN_3259 = imm_11_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire  imm_signBit_33 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_107 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_108 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_109 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_32 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_104 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_105 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_106 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_31 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_101 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_102 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_103 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_30 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_98 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_99 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_100 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_29 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_95 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_96 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_97 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_28 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_92 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_93 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_94 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_27 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_89 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_90 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_91 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [6:0] _imm_11_5_T_2 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _imm_11_5_T_1 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _imm_11_5_T = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _GEN_2461 = _T_447 ? inst[31:25] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [6:0] _GEN_2481 = _T_470 ? inst[31:25] : _GEN_2461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2501 = _T_494 ? inst[31:25] : _GEN_2481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] imm_11_5 = io_valid ? _GEN_2501 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [6:0] _GEN_3316 = imm_11_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [14:0] _T_497 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_498 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _imm_4_0_T_2 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_473 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_474 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _imm_4_0_T_1 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_450 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_451 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _imm_4_0_T = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_2465 = _T_447 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [4:0] _GEN_2485 = _T_470 ? inst[11:7] : _GEN_2465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2505 = _T_494 ? inst[11:7] : _GEN_2485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] imm_4_0 = io_valid ? _GEN_2505 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [4:0] _GEN_3317 = imm_4_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [11:0] _imm_T_85 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_26 = _imm_T_85[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_86 = imm_signBit_26; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_87 = imm_signBit_26 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_88 = {_imm_T_87,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [11:0] _imm_T_81 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_25 = _imm_T_85[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_82 = imm_signBit_26; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_83 = imm_signBit_26 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_84 = {_imm_T_87,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [11:0] _imm_T_77 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_24 = _imm_T_85[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_78 = imm_signBit_26; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_79 = imm_signBit_26 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_80 = {_imm_T_87,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_23 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_74 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_75 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_76 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_22 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_71 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_72 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_73 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_21 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_68 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_69 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_70 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_20 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_65 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_66 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_67 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_19 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_62 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_63 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_64 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _imm_12_T_5 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_4 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_3 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_2 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T_1 = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _imm_12_T = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _GEN_1789 = _T_182 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire  _GEN_1814 = _T_209 ? inst[31] : _GEN_1789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1839 = _T_236 ? inst[31] : _GEN_1814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1864 = _T_265 ? inst[31] : _GEN_1839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1889 = _T_292 ? inst[31] : _GEN_1864; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1914 = _T_321 ? inst[31] : _GEN_1889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_12 = io_valid & _GEN_1914; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire  _GEN_3309 = imm_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire [14:0] _T_325 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_326 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_327 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_6 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_296 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_297 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_298 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_5 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_269 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_270 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_271 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_4 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_240 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_241 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_242 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_3 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_213 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_214 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_215 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_2 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_186 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_187 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _T_188 = inst[7:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T_1 = inst[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_132 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_133 = 32'h6f == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [30:0] _T_134 = inst[30:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [20:0] _T_135 = inst[20:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _imm_11_T = inst[20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _GEN_1623 = _T_133 & inst[20]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire  _GEN_1795 = _T_182 ? inst[7] : _GEN_1623; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1820 = _T_209 ? inst[7] : _GEN_1795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1845 = _T_236 ? inst[7] : _GEN_1820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1870 = _T_265 ? inst[7] : _GEN_1845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1895 = _T_292 ? inst[7] : _GEN_1870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1920 = _T_321 ? inst[7] : _GEN_1895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_11 = io_valid & _GEN_1920; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire  _GEN_3302 = imm_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire [1:0] imm_hi_hi_6 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [5:0] _imm_10_5_T_5 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_4 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_3 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_2 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T_1 = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _imm_10_5_T = inst[30:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [5:0] _GEN_1790 = _T_182 ? inst[30:25] : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [5:0] _GEN_1815 = _T_209 ? inst[30:25] : _GEN_1790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1840 = _T_236 ? inst[30:25] : _GEN_1815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1865 = _T_265 ? inst[30:25] : _GEN_1840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1890 = _T_292 ? inst[30:25] : _GEN_1865; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1915 = _T_321 ? inst[30:25] : _GEN_1890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] imm_10_5 = io_valid ? _GEN_1915 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [5:0] _GEN_3310 = imm_10_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [7:0] imm_hi_6 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [3:0] _imm_4_1_T_5 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_4 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_3 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_2 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T_1 = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _imm_4_1_T = inst[11:8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [3:0] _GEN_1794 = _T_182 ? inst[11:8] : 4'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [3:0] _GEN_1819 = _T_209 ? inst[11:8] : _GEN_1794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1844 = _T_236 ? inst[11:8] : _GEN_1819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1869 = _T_265 ? inst[11:8] : _GEN_1844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1894 = _T_292 ? inst[11:8] : _GEN_1869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1919 = _T_321 ? inst[11:8] : _GEN_1894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] imm_4_1 = io_valid ? _GEN_1919 : 4'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [3:0] _GEN_3311 = imm_4_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [4:0] imm_lo_6 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_58 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_18 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_59 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_60 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_61 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_5 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_5 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_5 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_54 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_17 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_55 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_56 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_57 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_4 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_4 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_4 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_50 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_16 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_51 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_52 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_53 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_3 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_3 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_3 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_46 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_15 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_47 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_48 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_49 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_2 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_2 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_2 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_42 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_14 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_43 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_44 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_45 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [1:0] imm_hi_hi_1 = {imm_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [7:0] imm_hi_1 = {imm_12,imm_11,imm_10_5}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [4:0] imm_lo_1 = {imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire [12:0] _imm_T_38 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_13 = _imm_T_58[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_39 = imm_signBit_18; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [18:0] _imm_T_40 = imm_signBit_18 ? 19'h7ffff : 19'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_41 = {_imm_T_60,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_12 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_35 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_36 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_37 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _imm_20_T = inst[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire  _GEN_1621 = _T_133 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire  imm_20 = io_valid & _GEN_1621; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire  _GEN_3300 = imm_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire [19:0] _T_136 = inst[19:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [7:0] _imm_19_12_T = inst[19:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [7:0] _GEN_1624 = _T_133 ? inst[19:12] : 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [7:0] imm_19_12 = io_valid ? _GEN_1624 : 8'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [7:0] _GEN_3303 = imm_19_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [8:0] imm_hi_hi = {imm_20,imm_19_12}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire [9:0] imm_hi = {imm_20,imm_19_12,imm_11}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire [9:0] _imm_10_1_T = inst[30:21]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [9:0] _GEN_1622 = _T_133 ? inst[30:21] : 10'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [9:0] imm_10_1 = io_valid ? _GEN_1622 : 10'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [9:0] _GEN_3301 = imm_10_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [10:0] imm_lo = {imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire [20:0] _imm_T_31 = {imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire  imm_signBit_11 = _imm_T_31[20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_32 = imm_signBit_11; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [10:0] _imm_T_33 = imm_signBit_11 ? 11'h7ff : 11'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_34 = {_imm_T_33,imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _T_58 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_59 = 32'h17 == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _imm_31_12_T_1 = inst[31:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [31:0] _T_54 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_55 = 32'h37 == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _imm_31_12_T = inst[31:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [19:0] _GEN_704 = _T_55 ? inst[31:12] : 20'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [19:0] _GEN_773 = _T_59 ? inst[31:12] : _GEN_704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [19:0] imm_31_12 = io_valid ? _GEN_773 : 20'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [19:0] _GEN_3297 = imm_31_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [31:0] _imm_T_29 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire [31:0] _imm_T_30 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire [31:0] _imm_T_27 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire [31:0] _imm_T_28 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire  imm_signBit_8 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_24 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_25 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_26 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_7 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_21 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_22 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_23 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_6 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_18 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_19 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_20 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_5 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_15 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_16 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_17 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_4 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_12 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_13 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_14 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_3 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_9 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_10 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_11 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_2 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_6 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_7 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_8 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit_1 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T_3 = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_4 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_5 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  imm_signBit = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _imm_T = imm_signBit_33; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [19:0] _imm_T_1 = imm_signBit_33 ? 20'hfffff : 20'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _imm_T_2 = {_imm_T_108,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_70 = _T_1 ? _imm_T_109 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 22:24]
  wire [31:0] _GEN_141 = _T_7 ? _imm_T_109 : _GEN_70; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_212 = _T_13 ? _imm_T_109 : _GEN_141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_283 = _T_19 ? _imm_T_109 : _GEN_212; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_354 = _T_25 ? _imm_T_109 : _GEN_283; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_425 = _T_31 ? _imm_T_109 : _GEN_354; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_496 = _T_37 ? _imm_T_109 : _GEN_425; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_567 = _T_43 ? _imm_T_109 : _GEN_496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_638 = _T_49 ? _imm_T_109 : _GEN_567; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_707 = _T_55 ? _imm_T_29 : _GEN_638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [31:0] _GEN_776 = _T_59 ? _imm_T_29 : _GEN_707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [31:0] _GEN_1627 = _T_133 ? _imm_T_34 : _GEN_776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:127]
  wire [31:0] _GEN_1740 = _T_157 ? _imm_T_109 : _GEN_1627; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_1797 = _T_182 ? _imm_T_61 : _GEN_1740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1822 = _T_209 ? _imm_T_61 : _GEN_1797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1847 = _T_236 ? _imm_T_61 : _GEN_1822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1872 = _T_265 ? _imm_T_61 : _GEN_1847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1897 = _T_292 ? _imm_T_61 : _GEN_1872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_1922 = _T_321 ? _imm_T_61 : _GEN_1897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [31:0] _GEN_2003 = _T_348 ? _imm_T_109 : _GEN_1922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2116 = _T_368 ? _imm_T_109 : _GEN_2003; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2229 = _T_388 ? _imm_T_109 : _GEN_2116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2307 = _T_408 ? _imm_T_109 : _GEN_2229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2420 = _T_427 ? _imm_T_109 : _GEN_2307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2467 = _T_447 ? _imm_T_88 : _GEN_2420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [31:0] _GEN_2487 = _T_470 ? _imm_T_88 : _GEN_2467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [31:0] _GEN_2507 = _T_494 ? _imm_T_88 : _GEN_2487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [31:0] _GEN_2520 = _T_518 ? _imm_T_109 : _GEN_2507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2538 = _T_524 ? _imm_T_109 : _GEN_2520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_2549 = _T_533 ? _imm_T_109 : _GEN_2538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [31:0] _GEN_3135 = _T_595 ? _imm_T_109 : _GEN_2549; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_3156 = _T_602 ? _imm_T_109 : _GEN_3135; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _GEN_3170 = _T_609 ? _imm_T_109 : _GEN_3156; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28]
  wire [31:0] _GEN_3177 = _T_615 ? _imm_T_109 : _GEN_3170; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28]
  wire [31:0] imm = io_valid ? _GEN_3177 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [31:0] _GEN_3264 = imm; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [32:0] _T_432 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:47]
  wire [31:0] _T_433 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:47]
  wire [2:0] _T_438 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_439 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_442 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_436 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_437 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_440 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_434 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_435 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_441 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_443 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_445 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_423 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [4:0] _rs2_T_26 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_25 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_24 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_23 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_22 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_21 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_20 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_19 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_18 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_17 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_16 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_15 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_14 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_13 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_12 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_11 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_10 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_9 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_8 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_7 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_6 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_5 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_4 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_3 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_2 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T_1 = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _rs2_T = inst[24:20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_875 = _T_63 ? inst[24:20] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [4:0] _GEN_946 = _T_70 ? inst[24:20] : _GEN_875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1017 = _T_77 ? inst[24:20] : _GEN_946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1088 = _T_84 ? inst[24:20] : _GEN_1017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1159 = _T_91 ? inst[24:20] : _GEN_1088; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1230 = _T_98 ? inst[24:20] : _GEN_1159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1301 = _T_105 ? inst[24:20] : _GEN_1230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1372 = _T_112 ? inst[24:20] : _GEN_1301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1443 = _T_119 ? inst[24:20] : _GEN_1372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1514 = _T_126 ? inst[24:20] : _GEN_1443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1791 = _T_182 ? inst[24:20] : _GEN_1514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1816 = _T_209 ? inst[24:20] : _GEN_1791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1841 = _T_236 ? inst[24:20] : _GEN_1816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1866 = _T_265 ? inst[24:20] : _GEN_1841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1891 = _T_292 ? inst[24:20] : _GEN_1866; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1916 = _T_321 ? inst[24:20] : _GEN_1891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2462 = _T_447 ? inst[24:20] : _GEN_1916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2482 = _T_470 ? inst[24:20] : _GEN_2462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2502 = _T_494 ? inst[24:20] : _GEN_2482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2584 = _T_539 ? inst[24:20] : _GEN_2502; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2655 = _T_546 ? inst[24:20] : _GEN_2584; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2726 = _T_553 ? inst[24:20] : _GEN_2655; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2797 = _T_560 ? inst[24:20] : _GEN_2726; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2868 = _T_567 ? inst[24:20] : _GEN_2797; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2939 = _T_574 ? inst[24:20] : _GEN_2868; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3010 = _T_581 ? inst[24:20] : _GEN_2939; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3081 = _T_588 ? inst[24:20] : _GEN_3010; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs2 = io_valid ? _GEN_3081 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [4:0] _GEN_3299 = rs2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [2:0] _T_417 = rs2[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_418 = rs2[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_421 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_415 = rs2[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_416 = rs2[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_419 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_413 = rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_414 = ~rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_420 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_422 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_424 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_425 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 107:10]
  wire  _T_405 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_33 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_393 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:47]
  wire [31:0] _T_394 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:47]
  wire [2:0] _T_399 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_400 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_403 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_397 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_398 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_401 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_395 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_396 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_402 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_404 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_406 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_385 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_30 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_373 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:47]
  wire [31:0] _T_374 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:47]
  wire [2:0] _T_379 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_380 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_383 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_377 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_378 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_381 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_375 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_376 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_382 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_384 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_386 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_365 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_27 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_353 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:47]
  wire [31:0] _T_354 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:47]
  wire [2:0] _T_359 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_360 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_363 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_357 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_358 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_361 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_355 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_356 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_362 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_364 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_366 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _exceptionVec_WIRE_4 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_1995 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_2039 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2108 = _T_435 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2152 = _T_368 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2221 = _T_437 ? _GEN_2152 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2265 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2267 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2308 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2412 = _T_435 ? _GEN_2265 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2456 = _T_427 ? _GEN_2412 : _GEN_2265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  exceptionVec_4 = io_valid & _GEN_2456; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3315 = exceptionVec_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_4 = exceptionVec_4 ? 5'h4 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _T_512 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_44 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_500 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:47]
  wire [31:0] _T_501 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:47]
  wire [2:0] _T_506 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_507 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_510 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_504 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_505 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_508 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_502 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_503 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_509 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_511 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_513 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_488 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_41 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_476 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:47]
  wire [31:0] _T_477 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:47]
  wire [2:0] _T_482 = _T_433[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_483 = _T_433[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_486 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_480 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_481 = _T_433[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_484 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_478 = _T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_479 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_485 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_487 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_489 = ~_T_433[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_463 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [2:0] _T_457 = rs2[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_458 = rs2[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_461 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_455 = rs2[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_456 = rs2[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_459 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_453 = rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_454 = ~rs2[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_460 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_462 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_464 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_465 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 107:10]
  wire  _exceptionVec_WIRE_6 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2458 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 107:36 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_2468 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2478 = _T_435 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2492 = _T_470 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2498 = _T_437 ? _GEN_2492 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2512 = _T_494 ? _GEN_2498 : _GEN_2492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  exceptionVec_6 = io_valid & _GEN_2512; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3318 = exceptionVec_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_5 = exceptionVec_6 ? 5'h6 : _exceptionNO_T_4; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [1:0] now_internal_privilegeMode = io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_529 = 2'h3 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _exceptionVec_WIRE_8 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _T_530 = 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _T_531 = 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2523 = 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2527 = 2'h1 == io_now_internal_privilegeMode ? 1'h0 : 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2531 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : _GEN_2527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2542 = _T_524 & _GEN_2531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_8 = io_valid & _GEN_2542; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3326 = exceptionVec_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_6 = exceptionVec_8 ? 5'h8 : _exceptionNO_T_5; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_9 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2525 = 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2530 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2541 = _T_524 & _GEN_2530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_9 = io_valid & _GEN_2541; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3325 = exceptionVec_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_7 = exceptionVec_9 ? 5'h9 : _exceptionNO_T_6; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_11 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2528 = 2'h3 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2539 = _T_524 & _T_529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_11 = io_valid & _GEN_2539; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3324 = exceptionVec_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_8 = exceptionVec_11 ? 5'hb : _exceptionNO_T_7; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _now_reg_rs1_26 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _GEN_809 = io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_810 = 5'h1 == rs2 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_811 = 5'h2 == rs2 ? io_now_reg_2 : _GEN_810; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_812 = 5'h3 == rs2 ? io_now_reg_3 : _GEN_811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_813 = 5'h4 == rs2 ? io_now_reg_4 : _GEN_812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_814 = 5'h5 == rs2 ? io_now_reg_5 : _GEN_813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_815 = 5'h6 == rs2 ? io_now_reg_6 : _GEN_814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_816 = 5'h7 == rs2 ? io_now_reg_7 : _GEN_815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_817 = 5'h8 == rs2 ? io_now_reg_8 : _GEN_816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_818 = 5'h9 == rs2 ? io_now_reg_9 : _GEN_817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_819 = 5'ha == rs2 ? io_now_reg_10 : _GEN_818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_820 = 5'hb == rs2 ? io_now_reg_11 : _GEN_819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_821 = 5'hc == rs2 ? io_now_reg_12 : _GEN_820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_822 = 5'hd == rs2 ? io_now_reg_13 : _GEN_821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_823 = 5'he == rs2 ? io_now_reg_14 : _GEN_822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_824 = 5'hf == rs2 ? io_now_reg_15 : _GEN_823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_825 = 5'h10 == rs2 ? io_now_reg_16 : _GEN_824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_826 = 5'h11 == rs2 ? io_now_reg_17 : _GEN_825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_827 = 5'h12 == rs2 ? io_now_reg_18 : _GEN_826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_828 = 5'h13 == rs2 ? io_now_reg_19 : _GEN_827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_829 = 5'h14 == rs2 ? io_now_reg_20 : _GEN_828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_830 = 5'h15 == rs2 ? io_now_reg_21 : _GEN_829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_831 = 5'h16 == rs2 ? io_now_reg_22 : _GEN_830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_832 = 5'h17 == rs2 ? io_now_reg_23 : _GEN_831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_833 = 5'h18 == rs2 ? io_now_reg_24 : _GEN_832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_834 = 5'h19 == rs2 ? io_now_reg_25 : _GEN_833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_835 = 5'h1a == rs2 ? io_now_reg_26 : _GEN_834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_836 = 5'h1b == rs2 ? io_now_reg_27 : _GEN_835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_837 = 5'h1c == rs2 ? io_now_reg_28 : _GEN_836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_838 = 5'h1d == rs2 ? io_now_reg_29 : _GEN_837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_839 = 5'h1e == rs2 ? io_now_reg_30 : _GEN_838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _GEN_840 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _now_reg_rs2_14 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_329 = _GEN_31 >= _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:25]
  wire [31:0] now_csr_misa = io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_330 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_331 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_332 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_345 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] now_pc = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [32:0] _T_333 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:49]
  wire [31:0] _T_334 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:49]
  wire [2:0] _T_339 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_340 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_343 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_337 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_338 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_341 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_335 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_336 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_342 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_344 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_346 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_25 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _T_300 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:25]
  wire [31:0] _now_reg_rs2_13 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_301 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:48]
  wire  _T_302 = $signed(_T_300) >= $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:32]
  wire  _T_303 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_304 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_305 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_318 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_306 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:49]
  wire [31:0] _T_307 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:49]
  wire [2:0] _T_312 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_313 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_316 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_310 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_311 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_314 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_308 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_309 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_315 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_317 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_319 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_24 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_12 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_273 = _GEN_31 < _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:25]
  wire  _T_274 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_275 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_276 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_289 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_277 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:49]
  wire [31:0] _T_278 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:49]
  wire [2:0] _T_283 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_284 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_287 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_281 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_282 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_285 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_279 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_280 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_286 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_288 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_290 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_23 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _T_244 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:25]
  wire [31:0] _now_reg_rs2_11 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_245 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:47]
  wire  _T_246 = $signed(_T_300) < $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:32]
  wire  _T_247 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_248 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_249 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_262 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_250 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:49]
  wire [31:0] _T_251 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:49]
  wire [2:0] _T_256 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_257 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_260 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_254 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_255 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_258 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_252 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_253 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_259 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_261 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_263 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_22 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_10 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_217 = _GEN_31 != _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:25]
  wire  _T_218 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_219 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_220 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_233 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_221 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:49]
  wire [31:0] _T_222 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:49]
  wire [2:0] _T_227 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_228 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_231 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_225 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_226 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_229 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_223 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_224 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_230 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_232 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_234 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_21 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_9 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _T_190 = _GEN_31 == _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:25]
  wire  _T_191 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_192 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_193 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_206 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_194 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:49]
  wire [31:0] _T_195 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:49]
  wire [2:0] _T_200 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_201 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_204 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_198 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_199 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_202 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_196 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_197 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_203 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_205 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_207 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_162 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_163 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_164 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_179 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _now_reg_rs1_18 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_165 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:58]
  wire [31:0] _T_166 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:58]
  wire [30:0] _T_167 = _T_433[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:64]
  wire [31:0] _T_168 = {_T_433[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:43]
  wire [2:0] _T_173 = _T_168[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_174 = _T_168[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_177 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_171 = _T_168[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_172 = _T_168[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_175 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_169 = _T_168[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_170 = ~_T_168[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_176 = 2'h1 == _T_332 ? _T_170 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_178 = 2'h2 == _T_332 ? _T_172 : _T_176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_180 = 2'h3 == _T_332 ? _T_174 : _T_178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_139 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire  _T_140 = io_now_csr_misa[2]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:27]
  wire [1:0] _T_141 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire  _T_154 = 2'h3 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [32:0] _T_142 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:47]
  wire [31:0] _T_143 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:47]
  wire [2:0] _T_148 = _T_334[2:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:25]
  wire  _T_149 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_152 = 2'h2 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [1:0] _T_146 = _T_334[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:25]
  wire  _T_147 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_150 = 2'h1 == _T_332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_144 = _T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:25]
  wire  _T_145 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_151 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_153 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_155 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _exceptionVec_WIRE_0 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_1618 = _T_346 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_1663 = _T_133 & _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_1732 = _T_180 ? _GEN_1663 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1776 = _T_157 ? _GEN_1732 : _GEN_1663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1781 = _T_346 ? _GEN_1776 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1786 = _GEN_31 == _GEN_840 ? _GEN_1781 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1801 = _T_182 ? _GEN_1786 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1806 = _T_346 ? _GEN_1801 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1811 = _GEN_31 != _GEN_840 ? _GEN_1806 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1826 = _T_209 ? _GEN_1811 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1831 = _T_346 ? _GEN_1826 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1836 = $signed(_T_300) < $signed(_T_301) ? _GEN_1831 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1851 = _T_236 ? _GEN_1836 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1856 = _T_346 ? _GEN_1851 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1861 = _GEN_31 < _GEN_840 ? _GEN_1856 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1876 = _T_265 ? _GEN_1861 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1881 = _T_346 ? _GEN_1876 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1886 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1881 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1901 = _T_292 ? _GEN_1886 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1906 = _T_346 ? _GEN_1901 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1911 = _GEN_31 >= _GEN_840 ? _GEN_1906 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1926 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  exceptionVec_0 = io_valid & _GEN_1926; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3307 = exceptionVec_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_9 = exceptionVec_0 ? 5'h0 : _exceptionNO_T_8; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_64 = _T_1 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 125:24 128:24]
  wire  _GEN_135 = _T_7 ? 1'h0 : _GEN_64; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_206 = _T_13 ? 1'h0 : _GEN_135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_277 = _T_19 ? 1'h0 : _GEN_206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_348 = _T_25 ? 1'h0 : _GEN_277; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_419 = _T_31 ? 1'h0 : _GEN_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_490 = _T_37 ? 1'h0 : _GEN_419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_561 = _T_43 ? 1'h0 : _GEN_490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_632 = _T_49 ? 1'h0 : _GEN_561; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_703 = _T_55 ? 1'h0 : _GEN_632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_772 = _T_59 ? 1'h0 : _GEN_703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_873 = _T_63 ? 1'h0 : _GEN_772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_944 = _T_70 ? 1'h0 : _GEN_873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1015 = _T_77 ? 1'h0 : _GEN_944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1086 = _T_84 ? 1'h0 : _GEN_1015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1157 = _T_91 ? 1'h0 : _GEN_1086; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1228 = _T_98 ? 1'h0 : _GEN_1157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1299 = _T_105 ? 1'h0 : _GEN_1228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1370 = _T_112 ? 1'h0 : _GEN_1299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1441 = _T_119 ? 1'h0 : _GEN_1370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1512 = _T_126 ? 1'h0 : _GEN_1441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1620 = _T_133 ? 1'h0 : _GEN_1512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1734 = _T_157 ? 1'h0 : _GEN_1620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1788 = _T_182 ? 1'h0 : _GEN_1734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1813 = _T_209 ? 1'h0 : _GEN_1788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1838 = _T_236 ? 1'h0 : _GEN_1813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1863 = _T_265 ? 1'h0 : _GEN_1838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1888 = _T_292 ? 1'h0 : _GEN_1863; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1913 = _T_321 ? 1'h0 : _GEN_1888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1997 = _T_348 ? 1'h0 : _GEN_1913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2110 = _T_368 ? 1'h0 : _GEN_1997; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2223 = _T_388 ? 1'h0 : _GEN_2110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2301 = _T_408 ? 1'h0 : _GEN_2223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2414 = _T_427 ? 1'h0 : _GEN_2301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2460 = _T_447 ? 1'h0 : _GEN_2414; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2480 = _T_470 ? 1'h0 : _GEN_2460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2500 = _T_494 ? 1'h0 : _GEN_2480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2514 = _T_518 ? 1'h0 : _GEN_2500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2532 = _T_524 ? 1'h0 : _GEN_2514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2543 = _T_533 ? 1'h0 : _GEN_2532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2582 = _T_539 ? 1'h0 : _GEN_2543; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2653 = _T_546 ? 1'h0 : _GEN_2582; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2724 = _T_553 ? 1'h0 : _GEN_2653; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2795 = _T_560 ? 1'h0 : _GEN_2724; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2866 = _T_567 ? 1'h0 : _GEN_2795; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2937 = _T_574 ? 1'h0 : _GEN_2866; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3008 = _T_581 ? 1'h0 : _GEN_2937; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3079 = _T_588 ? 1'h0 : _GEN_3008; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3129 = _T_595 ? 1'h0 : _GEN_3079; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3150 = _T_602 ? 1'h0 : _GEN_3129; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3164 = _T_609 ? 1'h0 : _GEN_3150; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3171 = _T_615 ? 1'h0 : _GEN_3164; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  illegalInstruction = io_valid & _GEN_3171; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 119:36]
  wire  _GEN_3256 = illegalInstruction; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 119:36]
  wire  _T_607 = io_now_internal_privilegeMode == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:37]
  wire  illegalSret = io_now_internal_privilegeMode < 2'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 118:55]
  wire  _illegalSModeSret_T = io_now_internal_privilegeMode == 2'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 119:55]
  wire [31:0] now_csr_mstatus = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _mstatusOld_WIRE_1 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusOld_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_18 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _illegalSModeSret_T_1 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  illegalSModeSret = io_now_internal_privilegeMode == 2'h1 & mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 119:65]
  wire  _T_600 = illegalSret | illegalSModeSret; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:22]
  wire  _exceptionVec_WIRE_2 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_3118 = illegalSret | illegalSModeSret; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:22]
  wire  _GEN_3136 = _T_595 & _T_600; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3148 = io_now_internal_privilegeMode == 2'h3 ? _GEN_3136 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3162 = _T_602 ? _GEN_3148 : _GEN_3136; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_3179 = illegalInstruction | _GEN_3162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 144:33]
  wire  exceptionVec_2 = io_valid & _GEN_3179; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3327 = exceptionVec_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] _exceptionNO_T_10 = exceptionVec_2 ? 5'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_11 = exceptionVec_2 ? 5'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_12 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_12 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [4:0] _exceptionNO_T_12 = exceptionVec_2 ? 5'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _exceptionVec_WIRE_3 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _GEN_2521 = 32'h100073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  exceptionVec_3 = io_valid & _T_518; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3323 = exceptionVec_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [4:0] exceptionNO = exceptionVec_3 ? 5'h3 : _exceptionNO_T_10; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] now_csr_cycle = io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [32:0] _next_csr_cycle_T = io_now_csr_cycle + 32'h1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 126:37]
  wire [31:0] _next_csr_cycle_T_1 = io_now_csr_cycle + 32'h1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 126:37]
  wire [14:0] _T_3 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _funct3_T = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_4 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_5 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:63]
  wire [31:0] _next_reg_T_1 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:63]
  wire [14:0] _T_617 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_618 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_42 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_611 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_612 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_41 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_604 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_605 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_40 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_597 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_598 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_39 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_591 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_592 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_38 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_584 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_585 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_37 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_577 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_578 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_36 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_570 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_571 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_35 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_563 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_564 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_34 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_556 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_557 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_33 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_549 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_550 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_32 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_542 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_543 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_31 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_535 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_536 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_30 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_526 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_527 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_29 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_520 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_521 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_28 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_429 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_430 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_27 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_410 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_411 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_26 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_390 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_391 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_25 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_370 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_371 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_24 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_350 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_351 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_23 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_159 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_160 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_22 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_137 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_21 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_129 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_130 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_20 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_122 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_123 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_19 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_115 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_116 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_18 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_108 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_109 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_17 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_101 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_102 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_16 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_94 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_95 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_15 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_87 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_88 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_14 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_80 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_81 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_13 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_73 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_74 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_12 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_66 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_67 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_11 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_60 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_10 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [11:0] _T_56 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_9 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_51 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_52 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_8 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_45 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_46 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_7 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_39 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_40 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_6 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_33 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_34 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_5 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_27 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_28 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_4 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_21 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_22 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_3 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_15 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_16 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_2 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [14:0] _T_9 = inst[14:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [11:0] _T_10 = inst[11:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _rd_T_1 = inst[11:7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [4:0] _GEN_68 = _T_1 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [4:0] _GEN_139 = _T_7 ? inst[11:7] : _GEN_68; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_210 = _T_13 ? inst[11:7] : _GEN_139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_281 = _T_19 ? inst[11:7] : _GEN_210; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_352 = _T_25 ? inst[11:7] : _GEN_281; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_423 = _T_31 ? inst[11:7] : _GEN_352; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_494 = _T_37 ? inst[11:7] : _GEN_423; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_565 = _T_43 ? inst[11:7] : _GEN_494; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_636 = _T_49 ? inst[11:7] : _GEN_565; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_705 = _T_55 ? inst[11:7] : _GEN_636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_774 = _T_59 ? inst[11:7] : _GEN_705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_878 = _T_63 ? inst[11:7] : _GEN_774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_949 = _T_70 ? inst[11:7] : _GEN_878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1020 = _T_77 ? inst[11:7] : _GEN_949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1091 = _T_84 ? inst[11:7] : _GEN_1020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1162 = _T_91 ? inst[11:7] : _GEN_1091; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1233 = _T_98 ? inst[11:7] : _GEN_1162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1304 = _T_105 ? inst[11:7] : _GEN_1233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1375 = _T_112 ? inst[11:7] : _GEN_1304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1446 = _T_119 ? inst[11:7] : _GEN_1375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1517 = _T_126 ? inst[11:7] : _GEN_1446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1625 = _T_133 ? inst[11:7] : _GEN_1517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1738 = _T_157 ? inst[11:7] : _GEN_1625; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2001 = _T_348 ? inst[11:7] : _GEN_1738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2114 = _T_368 ? inst[11:7] : _GEN_2001; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2227 = _T_388 ? inst[11:7] : _GEN_2114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2305 = _T_408 ? inst[11:7] : _GEN_2227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2418 = _T_427 ? inst[11:7] : _GEN_2305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2518 = _T_518 ? inst[11:7] : _GEN_2418; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2536 = _T_524 ? inst[11:7] : _GEN_2518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2547 = _T_533 ? inst[11:7] : _GEN_2536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2587 = _T_539 ? inst[11:7] : _GEN_2547; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2658 = _T_546 ? inst[11:7] : _GEN_2587; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2729 = _T_553 ? inst[11:7] : _GEN_2658; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2800 = _T_560 ? inst[11:7] : _GEN_2729; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2871 = _T_567 ? inst[11:7] : _GEN_2800; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2942 = _T_574 ? inst[11:7] : _GEN_2871; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3013 = _T_581 ? inst[11:7] : _GEN_2942; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3084 = _T_588 ? inst[11:7] : _GEN_3013; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3133 = _T_595 ? inst[11:7] : _GEN_3084; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3154 = _T_602 ? inst[11:7] : _GEN_3133; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3168 = _T_609 ? inst[11:7] : _GEN_3154; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3175 = _T_615 ? inst[11:7] : _GEN_3168; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rd = io_valid ? _GEN_3175 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [4:0] _GEN_3262 = rd; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [31:0] _next_reg_rd = _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:63]
  wire [31:0] _GEN_32 = 5'h0 == rd ? _T_433 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_33 = 5'h1 == rd ? _T_433 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_34 = 5'h2 == rd ? _T_433 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_35 = 5'h3 == rd ? _T_433 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_36 = 5'h4 == rd ? _T_433 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_37 = 5'h5 == rd ? _T_433 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_38 = 5'h6 == rd ? _T_433 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_39 = 5'h7 == rd ? _T_433 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_40 = 5'h8 == rd ? _T_433 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_41 = 5'h9 == rd ? _T_433 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_42 = 5'ha == rd ? _T_433 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_43 = 5'hb == rd ? _T_433 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_44 = 5'hc == rd ? _T_433 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_45 = 5'hd == rd ? _T_433 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_46 = 5'he == rd ? _T_433 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_47 = 5'hf == rd ? _T_433 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_48 = 5'h10 == rd ? _T_433 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_49 = 5'h11 == rd ? _T_433 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_50 = 5'h12 == rd ? _T_433 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_51 = 5'h13 == rd ? _T_433 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_52 = 5'h14 == rd ? _T_433 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_53 = 5'h15 == rd ? _T_433 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_54 = 5'h16 == rd ? _T_433 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_55 = 5'h17 == rd ? _T_433 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_56 = 5'h18 == rd ? _T_433 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_57 = 5'h19 == rd ? _T_433 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_58 = 5'h1a == rd ? _T_433 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_59 = 5'h1b == rd ? _T_433 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_60 = 5'h1c == rd ? _T_433 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_61 = 5'h1d == rd ? _T_433 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_62 = 5'h1e == rd ? _T_433 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [31:0] _GEN_63 = 5'h1f == rd ? _T_433 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [2:0] _GEN_67 = _T_1 ? inst[14:12] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 18:24]
  wire [6:0] _GEN_69 = _T_1 ? inst[6:0] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 16:24]
  wire [31:0] _GEN_71 = _T_1 ? _GEN_32 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_72 = _T_1 ? _GEN_33 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_73 = _T_1 ? _GEN_34 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_74 = _T_1 ? _GEN_35 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_75 = _T_1 ? _GEN_36 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_76 = _T_1 ? _GEN_37 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_77 = _T_1 ? _GEN_38 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_78 = _T_1 ? _GEN_39 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_79 = _T_1 ? _GEN_40 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_80 = _T_1 ? _GEN_41 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_81 = _T_1 ? _GEN_42 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_82 = _T_1 ? _GEN_43 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_83 = _T_1 ? _GEN_44 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_84 = _T_1 ? _GEN_45 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_85 = _T_1 ? _GEN_46 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_86 = _T_1 ? _GEN_47 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_87 = _T_1 ? _GEN_48 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_88 = _T_1 ? _GEN_49 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_89 = _T_1 ? _GEN_50 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_90 = _T_1 ? _GEN_51 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_91 = _T_1 ? _GEN_52 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_92 = _T_1 ? _GEN_53 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_93 = _T_1 ? _GEN_54 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_94 = _T_1 ? _GEN_55 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_95 = _T_1 ? _GEN_56 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_96 = _T_1 ? _GEN_57 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_97 = _T_1 ? _GEN_58 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_98 = _T_1 ? _GEN_59 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_99 = _T_1 ? _GEN_60 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_100 = _T_1 ? _GEN_61 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_101 = _T_1 ? _GEN_62 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [31:0] _GEN_102 = _T_1 ? _GEN_63 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [2:0] _funct3_T_1 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_11 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_0 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_2 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:67]
  wire [31:0] _next_reg_T_3 = io_valid ? _GEN_3177 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:80]
  wire  _next_reg_T_4 = $signed(_T_300) < $signed(_next_reg_T_3); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:74]
  wire  _next_reg_T_5 = $signed(_T_300) < $signed(_next_reg_T_3); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:74]
  wire [31:0] _next_reg_rd_0 = {{31'd0}, $signed(_T_300) < $signed(_next_reg_T_3)}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_103 = 5'h0 == rd ? _next_reg_rd_0 : _GEN_71; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_104 = 5'h1 == rd ? _next_reg_rd_0 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_105 = 5'h2 == rd ? _next_reg_rd_0 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_106 = 5'h3 == rd ? _next_reg_rd_0 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_107 = 5'h4 == rd ? _next_reg_rd_0 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_108 = 5'h5 == rd ? _next_reg_rd_0 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_109 = 5'h6 == rd ? _next_reg_rd_0 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_110 = 5'h7 == rd ? _next_reg_rd_0 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_111 = 5'h8 == rd ? _next_reg_rd_0 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_112 = 5'h9 == rd ? _next_reg_rd_0 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_113 = 5'ha == rd ? _next_reg_rd_0 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_114 = 5'hb == rd ? _next_reg_rd_0 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_115 = 5'hc == rd ? _next_reg_rd_0 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_116 = 5'hd == rd ? _next_reg_rd_0 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_117 = 5'he == rd ? _next_reg_rd_0 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_118 = 5'hf == rd ? _next_reg_rd_0 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_119 = 5'h10 == rd ? _next_reg_rd_0 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_120 = 5'h11 == rd ? _next_reg_rd_0 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_121 = 5'h12 == rd ? _next_reg_rd_0 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_122 = 5'h13 == rd ? _next_reg_rd_0 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_123 = 5'h14 == rd ? _next_reg_rd_0 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_124 = 5'h15 == rd ? _next_reg_rd_0 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_125 = 5'h16 == rd ? _next_reg_rd_0 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_126 = 5'h17 == rd ? _next_reg_rd_0 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_127 = 5'h18 == rd ? _next_reg_rd_0 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_128 = 5'h19 == rd ? _next_reg_rd_0 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_129 = 5'h1a == rd ? _next_reg_rd_0 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_130 = 5'h1b == rd ? _next_reg_rd_0 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_131 = 5'h1c == rd ? _next_reg_rd_0 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_132 = 5'h1d == rd ? _next_reg_rd_0 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_133 = 5'h1e == rd ? _next_reg_rd_0 : _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [31:0] _GEN_134 = 5'h1f == rd ? _next_reg_rd_0 : _GEN_102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [2:0] _GEN_138 = _T_7 ? inst[14:12] : _GEN_67; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_140 = _T_7 ? inst[6:0] : _GEN_69; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_142 = _T_7 ? _GEN_103 : _GEN_71; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_143 = _T_7 ? _GEN_104 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_144 = _T_7 ? _GEN_105 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_145 = _T_7 ? _GEN_106 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_146 = _T_7 ? _GEN_107 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_147 = _T_7 ? _GEN_108 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_148 = _T_7 ? _GEN_109 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_149 = _T_7 ? _GEN_110 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_150 = _T_7 ? _GEN_111 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_151 = _T_7 ? _GEN_112 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_152 = _T_7 ? _GEN_113 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_153 = _T_7 ? _GEN_114 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_154 = _T_7 ? _GEN_115 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_155 = _T_7 ? _GEN_116 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_156 = _T_7 ? _GEN_117 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_157 = _T_7 ? _GEN_118 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_158 = _T_7 ? _GEN_119 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_159 = _T_7 ? _GEN_120 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_160 = _T_7 ? _GEN_121 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_161 = _T_7 ? _GEN_122 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_162 = _T_7 ? _GEN_123 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_163 = _T_7 ? _GEN_124 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_164 = _T_7 ? _GEN_125 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_165 = _T_7 ? _GEN_126 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_166 = _T_7 ? _GEN_127 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_167 = _T_7 ? _GEN_128 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_168 = _T_7 ? _GEN_129 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_169 = _T_7 ? _GEN_130 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_170 = _T_7 ? _GEN_131 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_171 = _T_7 ? _GEN_132 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_172 = _T_7 ? _GEN_133 : _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [31:0] _GEN_173 = _T_7 ? _GEN_134 : _GEN_102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [2:0] _funct3_T_2 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_17 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_1 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _next_reg_T_6 = _GEN_31 < imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:67]
  wire  _next_reg_T_7 = _GEN_31 < imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:67]
  wire [31:0] _next_reg_rd_1 = {{31'd0}, _GEN_31 < imm}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_174 = 5'h0 == rd ? _next_reg_rd_1 : _GEN_142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_175 = 5'h1 == rd ? _next_reg_rd_1 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_176 = 5'h2 == rd ? _next_reg_rd_1 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_177 = 5'h3 == rd ? _next_reg_rd_1 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_178 = 5'h4 == rd ? _next_reg_rd_1 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_179 = 5'h5 == rd ? _next_reg_rd_1 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_180 = 5'h6 == rd ? _next_reg_rd_1 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_181 = 5'h7 == rd ? _next_reg_rd_1 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_182 = 5'h8 == rd ? _next_reg_rd_1 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_183 = 5'h9 == rd ? _next_reg_rd_1 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_184 = 5'ha == rd ? _next_reg_rd_1 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_185 = 5'hb == rd ? _next_reg_rd_1 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_186 = 5'hc == rd ? _next_reg_rd_1 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_187 = 5'hd == rd ? _next_reg_rd_1 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_188 = 5'he == rd ? _next_reg_rd_1 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_189 = 5'hf == rd ? _next_reg_rd_1 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_190 = 5'h10 == rd ? _next_reg_rd_1 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_191 = 5'h11 == rd ? _next_reg_rd_1 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_192 = 5'h12 == rd ? _next_reg_rd_1 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_193 = 5'h13 == rd ? _next_reg_rd_1 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_194 = 5'h14 == rd ? _next_reg_rd_1 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_195 = 5'h15 == rd ? _next_reg_rd_1 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_196 = 5'h16 == rd ? _next_reg_rd_1 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_197 = 5'h17 == rd ? _next_reg_rd_1 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_198 = 5'h18 == rd ? _next_reg_rd_1 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_199 = 5'h19 == rd ? _next_reg_rd_1 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_200 = 5'h1a == rd ? _next_reg_rd_1 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_201 = 5'h1b == rd ? _next_reg_rd_1 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_202 = 5'h1c == rd ? _next_reg_rd_1 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_203 = 5'h1d == rd ? _next_reg_rd_1 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_204 = 5'h1e == rd ? _next_reg_rd_1 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [31:0] _GEN_205 = 5'h1f == rd ? _next_reg_rd_1 : _GEN_173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [2:0] _GEN_209 = _T_13 ? inst[14:12] : _GEN_138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_211 = _T_13 ? inst[6:0] : _GEN_140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_213 = _T_13 ? _GEN_174 : _GEN_142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_214 = _T_13 ? _GEN_175 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_215 = _T_13 ? _GEN_176 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_216 = _T_13 ? _GEN_177 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_217 = _T_13 ? _GEN_178 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_218 = _T_13 ? _GEN_179 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_219 = _T_13 ? _GEN_180 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_220 = _T_13 ? _GEN_181 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_221 = _T_13 ? _GEN_182 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_222 = _T_13 ? _GEN_183 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_223 = _T_13 ? _GEN_184 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_224 = _T_13 ? _GEN_185 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_225 = _T_13 ? _GEN_186 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_226 = _T_13 ? _GEN_187 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_227 = _T_13 ? _GEN_188 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_228 = _T_13 ? _GEN_189 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_229 = _T_13 ? _GEN_190 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_230 = _T_13 ? _GEN_191 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_231 = _T_13 ? _GEN_192 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_232 = _T_13 ? _GEN_193 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_233 = _T_13 ? _GEN_194 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_234 = _T_13 ? _GEN_195 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_235 = _T_13 ? _GEN_196 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_236 = _T_13 ? _GEN_197 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_237 = _T_13 ? _GEN_198 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_238 = _T_13 ? _GEN_199 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_239 = _T_13 ? _GEN_200 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_240 = _T_13 ? _GEN_201 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_241 = _T_13 ? _GEN_202 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_242 = _T_13 ? _GEN_203 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_243 = _T_13 ? _GEN_204 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [31:0] _GEN_244 = _T_13 ? _GEN_205 : _GEN_173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [2:0] _funct3_T_3 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_23 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_2 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_8 = _GEN_31 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:62]
  wire [31:0] _next_reg_rd_2 = _GEN_31 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:62]
  wire [31:0] _GEN_245 = 5'h0 == rd ? _next_reg_T_8 : _GEN_213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_246 = 5'h1 == rd ? _next_reg_T_8 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_247 = 5'h2 == rd ? _next_reg_T_8 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_248 = 5'h3 == rd ? _next_reg_T_8 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_249 = 5'h4 == rd ? _next_reg_T_8 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_250 = 5'h5 == rd ? _next_reg_T_8 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_251 = 5'h6 == rd ? _next_reg_T_8 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_252 = 5'h7 == rd ? _next_reg_T_8 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_253 = 5'h8 == rd ? _next_reg_T_8 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_254 = 5'h9 == rd ? _next_reg_T_8 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_255 = 5'ha == rd ? _next_reg_T_8 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_256 = 5'hb == rd ? _next_reg_T_8 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_257 = 5'hc == rd ? _next_reg_T_8 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_258 = 5'hd == rd ? _next_reg_T_8 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_259 = 5'he == rd ? _next_reg_T_8 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_260 = 5'hf == rd ? _next_reg_T_8 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_261 = 5'h10 == rd ? _next_reg_T_8 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_262 = 5'h11 == rd ? _next_reg_T_8 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_263 = 5'h12 == rd ? _next_reg_T_8 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_264 = 5'h13 == rd ? _next_reg_T_8 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_265 = 5'h14 == rd ? _next_reg_T_8 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_266 = 5'h15 == rd ? _next_reg_T_8 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_267 = 5'h16 == rd ? _next_reg_T_8 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_268 = 5'h17 == rd ? _next_reg_T_8 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_269 = 5'h18 == rd ? _next_reg_T_8 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_270 = 5'h19 == rd ? _next_reg_T_8 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_271 = 5'h1a == rd ? _next_reg_T_8 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_272 = 5'h1b == rd ? _next_reg_T_8 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_273 = 5'h1c == rd ? _next_reg_T_8 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_274 = 5'h1d == rd ? _next_reg_T_8 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_275 = 5'h1e == rd ? _next_reg_T_8 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [31:0] _GEN_276 = 5'h1f == rd ? _next_reg_T_8 : _GEN_244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [2:0] _GEN_280 = _T_19 ? inst[14:12] : _GEN_209; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_282 = _T_19 ? inst[6:0] : _GEN_211; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_284 = _T_19 ? _GEN_245 : _GEN_213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_285 = _T_19 ? _GEN_246 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_286 = _T_19 ? _GEN_247 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_287 = _T_19 ? _GEN_248 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_288 = _T_19 ? _GEN_249 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_289 = _T_19 ? _GEN_250 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_290 = _T_19 ? _GEN_251 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_291 = _T_19 ? _GEN_252 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_292 = _T_19 ? _GEN_253 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_293 = _T_19 ? _GEN_254 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_294 = _T_19 ? _GEN_255 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_295 = _T_19 ? _GEN_256 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_296 = _T_19 ? _GEN_257 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_297 = _T_19 ? _GEN_258 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_298 = _T_19 ? _GEN_259 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_299 = _T_19 ? _GEN_260 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_300 = _T_19 ? _GEN_261 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_301 = _T_19 ? _GEN_262 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_302 = _T_19 ? _GEN_263 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_303 = _T_19 ? _GEN_264 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_304 = _T_19 ? _GEN_265 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_305 = _T_19 ? _GEN_266 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_306 = _T_19 ? _GEN_267 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_307 = _T_19 ? _GEN_268 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_308 = _T_19 ? _GEN_269 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_309 = _T_19 ? _GEN_270 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_310 = _T_19 ? _GEN_271 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_311 = _T_19 ? _GEN_272 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_312 = _T_19 ? _GEN_273 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_313 = _T_19 ? _GEN_274 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_314 = _T_19 ? _GEN_275 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [31:0] _GEN_315 = _T_19 ? _GEN_276 : _GEN_244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [2:0] _funct3_T_4 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_29 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_3 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_9 = _GEN_31 | imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:62]
  wire [31:0] _next_reg_rd_3 = _GEN_31 | imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:62]
  wire [31:0] _GEN_316 = 5'h0 == rd ? _next_reg_T_9 : _GEN_284; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_317 = 5'h1 == rd ? _next_reg_T_9 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_318 = 5'h2 == rd ? _next_reg_T_9 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_319 = 5'h3 == rd ? _next_reg_T_9 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_320 = 5'h4 == rd ? _next_reg_T_9 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_321 = 5'h5 == rd ? _next_reg_T_9 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_322 = 5'h6 == rd ? _next_reg_T_9 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_323 = 5'h7 == rd ? _next_reg_T_9 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_324 = 5'h8 == rd ? _next_reg_T_9 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_325 = 5'h9 == rd ? _next_reg_T_9 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_326 = 5'ha == rd ? _next_reg_T_9 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_327 = 5'hb == rd ? _next_reg_T_9 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_328 = 5'hc == rd ? _next_reg_T_9 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_329 = 5'hd == rd ? _next_reg_T_9 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_330 = 5'he == rd ? _next_reg_T_9 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_331 = 5'hf == rd ? _next_reg_T_9 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_332 = 5'h10 == rd ? _next_reg_T_9 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_333 = 5'h11 == rd ? _next_reg_T_9 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_334 = 5'h12 == rd ? _next_reg_T_9 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_335 = 5'h13 == rd ? _next_reg_T_9 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_336 = 5'h14 == rd ? _next_reg_T_9 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_337 = 5'h15 == rd ? _next_reg_T_9 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_338 = 5'h16 == rd ? _next_reg_T_9 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_339 = 5'h17 == rd ? _next_reg_T_9 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_340 = 5'h18 == rd ? _next_reg_T_9 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_341 = 5'h19 == rd ? _next_reg_T_9 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_342 = 5'h1a == rd ? _next_reg_T_9 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_343 = 5'h1b == rd ? _next_reg_T_9 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_344 = 5'h1c == rd ? _next_reg_T_9 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_345 = 5'h1d == rd ? _next_reg_T_9 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_346 = 5'h1e == rd ? _next_reg_T_9 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [31:0] _GEN_347 = 5'h1f == rd ? _next_reg_T_9 : _GEN_315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [2:0] _GEN_351 = _T_25 ? inst[14:12] : _GEN_280; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_353 = _T_25 ? inst[6:0] : _GEN_282; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_355 = _T_25 ? _GEN_316 : _GEN_284; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_356 = _T_25 ? _GEN_317 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_357 = _T_25 ? _GEN_318 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_358 = _T_25 ? _GEN_319 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_359 = _T_25 ? _GEN_320 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_360 = _T_25 ? _GEN_321 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_361 = _T_25 ? _GEN_322 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_362 = _T_25 ? _GEN_323 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_363 = _T_25 ? _GEN_324 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_364 = _T_25 ? _GEN_325 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_365 = _T_25 ? _GEN_326 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_366 = _T_25 ? _GEN_327 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_367 = _T_25 ? _GEN_328 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_368 = _T_25 ? _GEN_329 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_369 = _T_25 ? _GEN_330 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_370 = _T_25 ? _GEN_331 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_371 = _T_25 ? _GEN_332 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_372 = _T_25 ? _GEN_333 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_373 = _T_25 ? _GEN_334 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_374 = _T_25 ? _GEN_335 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_375 = _T_25 ? _GEN_336 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_376 = _T_25 ? _GEN_337 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_377 = _T_25 ? _GEN_338 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_378 = _T_25 ? _GEN_339 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_379 = _T_25 ? _GEN_340 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_380 = _T_25 ? _GEN_341 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_381 = _T_25 ? _GEN_342 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_382 = _T_25 ? _GEN_343 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_383 = _T_25 ? _GEN_344 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_384 = _T_25 ? _GEN_345 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_385 = _T_25 ? _GEN_346 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [31:0] _GEN_386 = _T_25 ? _GEN_347 : _GEN_315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [2:0] _funct3_T_5 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_35 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_4 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_10 = _GEN_31 ^ imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:62]
  wire [31:0] _next_reg_rd_4 = _GEN_31 ^ imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:62]
  wire [31:0] _GEN_387 = 5'h0 == rd ? _next_reg_T_10 : _GEN_355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_388 = 5'h1 == rd ? _next_reg_T_10 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_389 = 5'h2 == rd ? _next_reg_T_10 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_390 = 5'h3 == rd ? _next_reg_T_10 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_391 = 5'h4 == rd ? _next_reg_T_10 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_392 = 5'h5 == rd ? _next_reg_T_10 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_393 = 5'h6 == rd ? _next_reg_T_10 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_394 = 5'h7 == rd ? _next_reg_T_10 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_395 = 5'h8 == rd ? _next_reg_T_10 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_396 = 5'h9 == rd ? _next_reg_T_10 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_397 = 5'ha == rd ? _next_reg_T_10 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_398 = 5'hb == rd ? _next_reg_T_10 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_399 = 5'hc == rd ? _next_reg_T_10 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_400 = 5'hd == rd ? _next_reg_T_10 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_401 = 5'he == rd ? _next_reg_T_10 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_402 = 5'hf == rd ? _next_reg_T_10 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_403 = 5'h10 == rd ? _next_reg_T_10 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_404 = 5'h11 == rd ? _next_reg_T_10 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_405 = 5'h12 == rd ? _next_reg_T_10 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_406 = 5'h13 == rd ? _next_reg_T_10 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_407 = 5'h14 == rd ? _next_reg_T_10 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_408 = 5'h15 == rd ? _next_reg_T_10 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_409 = 5'h16 == rd ? _next_reg_T_10 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_410 = 5'h17 == rd ? _next_reg_T_10 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_411 = 5'h18 == rd ? _next_reg_T_10 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_412 = 5'h19 == rd ? _next_reg_T_10 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_413 = 5'h1a == rd ? _next_reg_T_10 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_414 = 5'h1b == rd ? _next_reg_T_10 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_415 = 5'h1c == rd ? _next_reg_T_10 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_416 = 5'h1d == rd ? _next_reg_T_10 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_417 = 5'h1e == rd ? _next_reg_T_10 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [31:0] _GEN_418 = 5'h1f == rd ? _next_reg_T_10 : _GEN_386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [2:0] _GEN_422 = _T_31 ? inst[14:12] : _GEN_351; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_424 = _T_31 ? inst[6:0] : _GEN_353; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_426 = _T_31 ? _GEN_387 : _GEN_355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_427 = _T_31 ? _GEN_388 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_428 = _T_31 ? _GEN_389 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_429 = _T_31 ? _GEN_390 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_430 = _T_31 ? _GEN_391 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_431 = _T_31 ? _GEN_392 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_432 = _T_31 ? _GEN_393 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_433 = _T_31 ? _GEN_394 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_434 = _T_31 ? _GEN_395 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_435 = _T_31 ? _GEN_396 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_436 = _T_31 ? _GEN_397 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_437 = _T_31 ? _GEN_398 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_438 = _T_31 ? _GEN_399 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_439 = _T_31 ? _GEN_400 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_440 = _T_31 ? _GEN_401 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_441 = _T_31 ? _GEN_402 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_442 = _T_31 ? _GEN_403 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_443 = _T_31 ? _GEN_404 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_444 = _T_31 ? _GEN_405 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_445 = _T_31 ? _GEN_406 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_446 = _T_31 ? _GEN_407 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_447 = _T_31 ? _GEN_408 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_448 = _T_31 ? _GEN_409 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_449 = _T_31 ? _GEN_410 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_450 = _T_31 ? _GEN_411 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_451 = _T_31 ? _GEN_412 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_452 = _T_31 ? _GEN_413 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_453 = _T_31 ? _GEN_414 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_454 = _T_31 ? _GEN_415 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_455 = _T_31 ? _GEN_416 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_456 = _T_31 ? _GEN_417 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [31:0] _GEN_457 = _T_31 ? _GEN_418 : _GEN_386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [2:0] _funct3_T_6 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_41 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _next_reg_T_11 = imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:68]
  wire [31:0] _now_reg_rs1_5 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [62:0] _GEN_3347 = {{31'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [62:0] _next_reg_T_12 = _GEN_3347 << imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [31:0] _next_reg_rd_5 = _next_reg_T_12[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_458 = 5'h0 == rd ? _next_reg_T_12[31:0] : _GEN_426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_459 = 5'h1 == rd ? _next_reg_T_12[31:0] : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_460 = 5'h2 == rd ? _next_reg_T_12[31:0] : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_461 = 5'h3 == rd ? _next_reg_T_12[31:0] : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_462 = 5'h4 == rd ? _next_reg_T_12[31:0] : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_463 = 5'h5 == rd ? _next_reg_T_12[31:0] : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_464 = 5'h6 == rd ? _next_reg_T_12[31:0] : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_465 = 5'h7 == rd ? _next_reg_T_12[31:0] : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_466 = 5'h8 == rd ? _next_reg_T_12[31:0] : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_467 = 5'h9 == rd ? _next_reg_T_12[31:0] : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_468 = 5'ha == rd ? _next_reg_T_12[31:0] : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_469 = 5'hb == rd ? _next_reg_T_12[31:0] : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_470 = 5'hc == rd ? _next_reg_T_12[31:0] : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_471 = 5'hd == rd ? _next_reg_T_12[31:0] : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_472 = 5'he == rd ? _next_reg_T_12[31:0] : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_473 = 5'hf == rd ? _next_reg_T_12[31:0] : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_474 = 5'h10 == rd ? _next_reg_T_12[31:0] : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_475 = 5'h11 == rd ? _next_reg_T_12[31:0] : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_476 = 5'h12 == rd ? _next_reg_T_12[31:0] : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_477 = 5'h13 == rd ? _next_reg_T_12[31:0] : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_478 = 5'h14 == rd ? _next_reg_T_12[31:0] : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_479 = 5'h15 == rd ? _next_reg_T_12[31:0] : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_480 = 5'h16 == rd ? _next_reg_T_12[31:0] : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_481 = 5'h17 == rd ? _next_reg_T_12[31:0] : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_482 = 5'h18 == rd ? _next_reg_T_12[31:0] : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_483 = 5'h19 == rd ? _next_reg_T_12[31:0] : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_484 = 5'h1a == rd ? _next_reg_T_12[31:0] : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_485 = 5'h1b == rd ? _next_reg_T_12[31:0] : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_486 = 5'h1c == rd ? _next_reg_T_12[31:0] : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_487 = 5'h1d == rd ? _next_reg_T_12[31:0] : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_488 = 5'h1e == rd ? _next_reg_T_12[31:0] : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [31:0] _GEN_489 = 5'h1f == rd ? _next_reg_T_12[31:0] : _GEN_457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [2:0] _GEN_493 = _T_37 ? inst[14:12] : _GEN_422; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_495 = _T_37 ? inst[6:0] : _GEN_424; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_497 = _T_37 ? _GEN_458 : _GEN_426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_498 = _T_37 ? _GEN_459 : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_499 = _T_37 ? _GEN_460 : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_500 = _T_37 ? _GEN_461 : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_501 = _T_37 ? _GEN_462 : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_502 = _T_37 ? _GEN_463 : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_503 = _T_37 ? _GEN_464 : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_504 = _T_37 ? _GEN_465 : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_505 = _T_37 ? _GEN_466 : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_506 = _T_37 ? _GEN_467 : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_507 = _T_37 ? _GEN_468 : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_508 = _T_37 ? _GEN_469 : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_509 = _T_37 ? _GEN_470 : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_510 = _T_37 ? _GEN_471 : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_511 = _T_37 ? _GEN_472 : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_512 = _T_37 ? _GEN_473 : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_513 = _T_37 ? _GEN_474 : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_514 = _T_37 ? _GEN_475 : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_515 = _T_37 ? _GEN_476 : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_516 = _T_37 ? _GEN_477 : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_517 = _T_37 ? _GEN_478 : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_518 = _T_37 ? _GEN_479 : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_519 = _T_37 ? _GEN_480 : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_520 = _T_37 ? _GEN_481 : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_521 = _T_37 ? _GEN_482 : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_522 = _T_37 ? _GEN_483 : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_523 = _T_37 ? _GEN_484 : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_524 = _T_37 ? _GEN_485 : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_525 = _T_37 ? _GEN_486 : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_526 = _T_37 ? _GEN_487 : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_527 = _T_37 ? _GEN_488 : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [31:0] _GEN_528 = _T_37 ? _GEN_489 : _GEN_457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [2:0] _funct3_T_7 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_47 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [4:0] _next_reg_T_13 = imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:68]
  wire [31:0] _now_reg_rs1_6 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_14 = _GEN_31 >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:62]
  wire [31:0] _next_reg_rd_6 = _GEN_31 >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:62]
  wire [31:0] _GEN_529 = 5'h0 == rd ? _next_reg_T_14 : _GEN_497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_530 = 5'h1 == rd ? _next_reg_T_14 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_531 = 5'h2 == rd ? _next_reg_T_14 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_532 = 5'h3 == rd ? _next_reg_T_14 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_533 = 5'h4 == rd ? _next_reg_T_14 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_534 = 5'h5 == rd ? _next_reg_T_14 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_535 = 5'h6 == rd ? _next_reg_T_14 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_536 = 5'h7 == rd ? _next_reg_T_14 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_537 = 5'h8 == rd ? _next_reg_T_14 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_538 = 5'h9 == rd ? _next_reg_T_14 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_539 = 5'ha == rd ? _next_reg_T_14 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_540 = 5'hb == rd ? _next_reg_T_14 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_541 = 5'hc == rd ? _next_reg_T_14 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_542 = 5'hd == rd ? _next_reg_T_14 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_543 = 5'he == rd ? _next_reg_T_14 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_544 = 5'hf == rd ? _next_reg_T_14 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_545 = 5'h10 == rd ? _next_reg_T_14 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_546 = 5'h11 == rd ? _next_reg_T_14 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_547 = 5'h12 == rd ? _next_reg_T_14 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_548 = 5'h13 == rd ? _next_reg_T_14 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_549 = 5'h14 == rd ? _next_reg_T_14 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_550 = 5'h15 == rd ? _next_reg_T_14 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_551 = 5'h16 == rd ? _next_reg_T_14 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_552 = 5'h17 == rd ? _next_reg_T_14 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_553 = 5'h18 == rd ? _next_reg_T_14 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_554 = 5'h19 == rd ? _next_reg_T_14 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_555 = 5'h1a == rd ? _next_reg_T_14 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_556 = 5'h1b == rd ? _next_reg_T_14 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_557 = 5'h1c == rd ? _next_reg_T_14 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_558 = 5'h1d == rd ? _next_reg_T_14 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_559 = 5'h1e == rd ? _next_reg_T_14 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [31:0] _GEN_560 = 5'h1f == rd ? _next_reg_T_14 : _GEN_528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [2:0] _GEN_564 = _T_43 ? inst[14:12] : _GEN_493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_566 = _T_43 ? inst[6:0] : _GEN_495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_568 = _T_43 ? _GEN_529 : _GEN_497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_569 = _T_43 ? _GEN_530 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_570 = _T_43 ? _GEN_531 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_571 = _T_43 ? _GEN_532 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_572 = _T_43 ? _GEN_533 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_573 = _T_43 ? _GEN_534 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_574 = _T_43 ? _GEN_535 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_575 = _T_43 ? _GEN_536 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_576 = _T_43 ? _GEN_537 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_577 = _T_43 ? _GEN_538 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_578 = _T_43 ? _GEN_539 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_579 = _T_43 ? _GEN_540 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_580 = _T_43 ? _GEN_541 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_581 = _T_43 ? _GEN_542 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_582 = _T_43 ? _GEN_543 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_583 = _T_43 ? _GEN_544 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_584 = _T_43 ? _GEN_545 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_585 = _T_43 ? _GEN_546 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_586 = _T_43 ? _GEN_547 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_587 = _T_43 ? _GEN_548 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_588 = _T_43 ? _GEN_549 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_589 = _T_43 ? _GEN_550 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_590 = _T_43 ? _GEN_551 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_591 = _T_43 ? _GEN_552 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_592 = _T_43 ? _GEN_553 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_593 = _T_43 ? _GEN_554 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_594 = _T_43 ? _GEN_555 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_595 = _T_43 ? _GEN_556 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_596 = _T_43 ? _GEN_557 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_597 = _T_43 ? _GEN_558 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_598 = _T_43 ? _GEN_559 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [31:0] _GEN_599 = _T_43 ? _GEN_560 : _GEN_528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [2:0] _funct3_T_8 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_53 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_7 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_15 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:63]
  wire [4:0] _next_reg_T_16 = imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:76]
  wire [31:0] _next_reg_T_17 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:70]
  wire [31:0] _next_reg_T_18 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:84]
  wire [31:0] _next_reg_rd_7 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:84]
  wire [31:0] _GEN_600 = 5'h0 == rd ? _next_reg_T_18 : _GEN_568; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_601 = 5'h1 == rd ? _next_reg_T_18 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_602 = 5'h2 == rd ? _next_reg_T_18 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_603 = 5'h3 == rd ? _next_reg_T_18 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_604 = 5'h4 == rd ? _next_reg_T_18 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_605 = 5'h5 == rd ? _next_reg_T_18 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_606 = 5'h6 == rd ? _next_reg_T_18 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_607 = 5'h7 == rd ? _next_reg_T_18 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_608 = 5'h8 == rd ? _next_reg_T_18 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_609 = 5'h9 == rd ? _next_reg_T_18 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_610 = 5'ha == rd ? _next_reg_T_18 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_611 = 5'hb == rd ? _next_reg_T_18 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_612 = 5'hc == rd ? _next_reg_T_18 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_613 = 5'hd == rd ? _next_reg_T_18 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_614 = 5'he == rd ? _next_reg_T_18 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_615 = 5'hf == rd ? _next_reg_T_18 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_616 = 5'h10 == rd ? _next_reg_T_18 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_617 = 5'h11 == rd ? _next_reg_T_18 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_618 = 5'h12 == rd ? _next_reg_T_18 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_619 = 5'h13 == rd ? _next_reg_T_18 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_620 = 5'h14 == rd ? _next_reg_T_18 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_621 = 5'h15 == rd ? _next_reg_T_18 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_622 = 5'h16 == rd ? _next_reg_T_18 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_623 = 5'h17 == rd ? _next_reg_T_18 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_624 = 5'h18 == rd ? _next_reg_T_18 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_625 = 5'h19 == rd ? _next_reg_T_18 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_626 = 5'h1a == rd ? _next_reg_T_18 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_627 = 5'h1b == rd ? _next_reg_T_18 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_628 = 5'h1c == rd ? _next_reg_T_18 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_629 = 5'h1d == rd ? _next_reg_T_18 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_630 = 5'h1e == rd ? _next_reg_T_18 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [31:0] _GEN_631 = 5'h1f == rd ? _next_reg_T_18 : _GEN_599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [2:0] _GEN_635 = _T_49 ? inst[14:12] : _GEN_564; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_637 = _T_49 ? inst[6:0] : _GEN_566; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_639 = _T_49 ? _GEN_600 : _GEN_568; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_640 = _T_49 ? _GEN_601 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_641 = _T_49 ? _GEN_602 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_642 = _T_49 ? _GEN_603 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_643 = _T_49 ? _GEN_604 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_644 = _T_49 ? _GEN_605 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_645 = _T_49 ? _GEN_606 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_646 = _T_49 ? _GEN_607 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_647 = _T_49 ? _GEN_608 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_648 = _T_49 ? _GEN_609 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_649 = _T_49 ? _GEN_610 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_650 = _T_49 ? _GEN_611 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_651 = _T_49 ? _GEN_612 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_652 = _T_49 ? _GEN_613 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_653 = _T_49 ? _GEN_614 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_654 = _T_49 ? _GEN_615 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_655 = _T_49 ? _GEN_616 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_656 = _T_49 ? _GEN_617 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_657 = _T_49 ? _GEN_618 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_658 = _T_49 ? _GEN_619 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_659 = _T_49 ? _GEN_620 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_660 = _T_49 ? _GEN_621 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_661 = _T_49 ? _GEN_622 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_662 = _T_49 ? _GEN_623 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_663 = _T_49 ? _GEN_624 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_664 = _T_49 ? _GEN_625 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_665 = _T_49 ? _GEN_626 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_666 = _T_49 ? _GEN_627 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_667 = _T_49 ? _GEN_628 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_668 = _T_49 ? _GEN_629 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_669 = _T_49 ? _GEN_630 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [31:0] _GEN_670 = _T_49 ? _GEN_631 : _GEN_599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [6:0] _T_57 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  imm_signBit_9 = _imm_T_29[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_rd_8 = imm; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [31:0] _GEN_671 = 5'h0 == rd ? imm : _GEN_639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_672 = 5'h1 == rd ? imm : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_673 = 5'h2 == rd ? imm : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_674 = 5'h3 == rd ? imm : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_675 = 5'h4 == rd ? imm : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_676 = 5'h5 == rd ? imm : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_677 = 5'h6 == rd ? imm : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_678 = 5'h7 == rd ? imm : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_679 = 5'h8 == rd ? imm : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_680 = 5'h9 == rd ? imm : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_681 = 5'ha == rd ? imm : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_682 = 5'hb == rd ? imm : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_683 = 5'hc == rd ? imm : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_684 = 5'hd == rd ? imm : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_685 = 5'he == rd ? imm : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_686 = 5'hf == rd ? imm : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_687 = 5'h10 == rd ? imm : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_688 = 5'h11 == rd ? imm : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_689 = 5'h12 == rd ? imm : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_690 = 5'h13 == rd ? imm : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_691 = 5'h14 == rd ? imm : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_692 = 5'h15 == rd ? imm : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_693 = 5'h16 == rd ? imm : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_694 = 5'h17 == rd ? imm : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_695 = 5'h18 == rd ? imm : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_696 = 5'h19 == rd ? imm : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_697 = 5'h1a == rd ? imm : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_698 = 5'h1b == rd ? imm : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_699 = 5'h1c == rd ? imm : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_700 = 5'h1d == rd ? imm : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_701 = 5'h1e == rd ? imm : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [31:0] _GEN_702 = 5'h1f == rd ? imm : _GEN_670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [6:0] _GEN_706 = _T_55 ? inst[6:0] : _GEN_637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_708 = _T_55 ? _GEN_671 : _GEN_639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_709 = _T_55 ? _GEN_672 : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_710 = _T_55 ? _GEN_673 : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_711 = _T_55 ? _GEN_674 : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_712 = _T_55 ? _GEN_675 : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_713 = _T_55 ? _GEN_676 : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_714 = _T_55 ? _GEN_677 : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_715 = _T_55 ? _GEN_678 : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_716 = _T_55 ? _GEN_679 : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_717 = _T_55 ? _GEN_680 : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_718 = _T_55 ? _GEN_681 : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_719 = _T_55 ? _GEN_682 : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_720 = _T_55 ? _GEN_683 : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_721 = _T_55 ? _GEN_684 : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_722 = _T_55 ? _GEN_685 : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_723 = _T_55 ? _GEN_686 : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_724 = _T_55 ? _GEN_687 : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_725 = _T_55 ? _GEN_688 : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_726 = _T_55 ? _GEN_689 : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_727 = _T_55 ? _GEN_690 : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_728 = _T_55 ? _GEN_691 : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_729 = _T_55 ? _GEN_692 : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_730 = _T_55 ? _GEN_693 : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_731 = _T_55 ? _GEN_694 : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_732 = _T_55 ? _GEN_695 : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_733 = _T_55 ? _GEN_696 : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_734 = _T_55 ? _GEN_697 : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_735 = _T_55 ? _GEN_698 : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_736 = _T_55 ? _GEN_699 : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_737 = _T_55 ? _GEN_700 : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_738 = _T_55 ? _GEN_701 : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [31:0] _GEN_739 = _T_55 ? _GEN_702 : _GEN_670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [6:0] _T_61 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  imm_signBit_10 = _imm_T_29[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [32:0] _next_reg_T_19 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:57]
  wire [31:0] _next_reg_T_20 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:57]
  wire [31:0] _next_reg_rd_9 = _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:57]
  wire [31:0] _GEN_740 = 5'h0 == rd ? _T_334 : _GEN_708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_741 = 5'h1 == rd ? _T_334 : _GEN_709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_742 = 5'h2 == rd ? _T_334 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_743 = 5'h3 == rd ? _T_334 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_744 = 5'h4 == rd ? _T_334 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_745 = 5'h5 == rd ? _T_334 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_746 = 5'h6 == rd ? _T_334 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_747 = 5'h7 == rd ? _T_334 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_748 = 5'h8 == rd ? _T_334 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_749 = 5'h9 == rd ? _T_334 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_750 = 5'ha == rd ? _T_334 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_751 = 5'hb == rd ? _T_334 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_752 = 5'hc == rd ? _T_334 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_753 = 5'hd == rd ? _T_334 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_754 = 5'he == rd ? _T_334 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_755 = 5'hf == rd ? _T_334 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_756 = 5'h10 == rd ? _T_334 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_757 = 5'h11 == rd ? _T_334 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_758 = 5'h12 == rd ? _T_334 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_759 = 5'h13 == rd ? _T_334 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_760 = 5'h14 == rd ? _T_334 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_761 = 5'h15 == rd ? _T_334 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_762 = 5'h16 == rd ? _T_334 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_763 = 5'h17 == rd ? _T_334 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_764 = 5'h18 == rd ? _T_334 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_765 = 5'h19 == rd ? _T_334 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_766 = 5'h1a == rd ? _T_334 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_767 = 5'h1b == rd ? _T_334 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_768 = 5'h1c == rd ? _T_334 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_769 = 5'h1d == rd ? _T_334 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_770 = 5'h1e == rd ? _T_334 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [31:0] _GEN_771 = 5'h1f == rd ? _T_334 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [6:0] _GEN_775 = _T_59 ? inst[6:0] : _GEN_706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_777 = _T_59 ? _GEN_740 : _GEN_708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_778 = _T_59 ? _GEN_741 : _GEN_709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_779 = _T_59 ? _GEN_742 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_780 = _T_59 ? _GEN_743 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_781 = _T_59 ? _GEN_744 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_782 = _T_59 ? _GEN_745 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_783 = _T_59 ? _GEN_746 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_784 = _T_59 ? _GEN_747 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_785 = _T_59 ? _GEN_748 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_786 = _T_59 ? _GEN_749 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_787 = _T_59 ? _GEN_750 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_788 = _T_59 ? _GEN_751 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_789 = _T_59 ? _GEN_752 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_790 = _T_59 ? _GEN_753 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_791 = _T_59 ? _GEN_754 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_792 = _T_59 ? _GEN_755 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_793 = _T_59 ? _GEN_756 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_794 = _T_59 ? _GEN_757 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_795 = _T_59 ? _GEN_758 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_796 = _T_59 ? _GEN_759 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_797 = _T_59 ? _GEN_760 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_798 = _T_59 ? _GEN_761 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_799 = _T_59 ? _GEN_762 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_800 = _T_59 ? _GEN_763 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_801 = _T_59 ? _GEN_764 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_802 = _T_59 ? _GEN_765 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_803 = _T_59 ? _GEN_766 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_804 = _T_59 ? _GEN_767 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_805 = _T_59 ? _GEN_768 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_806 = _T_59 ? _GEN_769 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_807 = _T_59 ? _GEN_770 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [31:0] _GEN_808 = _T_59 ? _GEN_771 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [6:0] _funct7_T = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_9 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_68 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_8 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_21 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [31:0] _next_reg_T_22 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [31:0] _next_reg_rd_10 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [31:0] _GEN_841 = 5'h0 == rd ? _next_reg_T_22 : _GEN_777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_842 = 5'h1 == rd ? _next_reg_T_22 : _GEN_778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_843 = 5'h2 == rd ? _next_reg_T_22 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_844 = 5'h3 == rd ? _next_reg_T_22 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_845 = 5'h4 == rd ? _next_reg_T_22 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_846 = 5'h5 == rd ? _next_reg_T_22 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_847 = 5'h6 == rd ? _next_reg_T_22 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_848 = 5'h7 == rd ? _next_reg_T_22 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_849 = 5'h8 == rd ? _next_reg_T_22 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_850 = 5'h9 == rd ? _next_reg_T_22 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_851 = 5'ha == rd ? _next_reg_T_22 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_852 = 5'hb == rd ? _next_reg_T_22 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_853 = 5'hc == rd ? _next_reg_T_22 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_854 = 5'hd == rd ? _next_reg_T_22 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_855 = 5'he == rd ? _next_reg_T_22 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_856 = 5'hf == rd ? _next_reg_T_22 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_857 = 5'h10 == rd ? _next_reg_T_22 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_858 = 5'h11 == rd ? _next_reg_T_22 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_859 = 5'h12 == rd ? _next_reg_T_22 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_860 = 5'h13 == rd ? _next_reg_T_22 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_861 = 5'h14 == rd ? _next_reg_T_22 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_862 = 5'h15 == rd ? _next_reg_T_22 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_863 = 5'h16 == rd ? _next_reg_T_22 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_864 = 5'h17 == rd ? _next_reg_T_22 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_865 = 5'h18 == rd ? _next_reg_T_22 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_866 = 5'h19 == rd ? _next_reg_T_22 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_867 = 5'h1a == rd ? _next_reg_T_22 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_868 = 5'h1b == rd ? _next_reg_T_22 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_869 = 5'h1c == rd ? _next_reg_T_22 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_870 = 5'h1d == rd ? _next_reg_T_22 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_871 = 5'h1e == rd ? _next_reg_T_22 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [31:0] _GEN_872 = 5'h1f == rd ? _next_reg_T_22 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [6:0] _GEN_874 = _T_63 ? inst[31:25] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 21:24]
  wire [2:0] _GEN_877 = _T_63 ? inst[14:12] : _GEN_635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_879 = _T_63 ? inst[6:0] : _GEN_775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_880 = _T_63 ? _GEN_841 : _GEN_777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_881 = _T_63 ? _GEN_842 : _GEN_778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_882 = _T_63 ? _GEN_843 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_883 = _T_63 ? _GEN_844 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_884 = _T_63 ? _GEN_845 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_885 = _T_63 ? _GEN_846 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_886 = _T_63 ? _GEN_847 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_887 = _T_63 ? _GEN_848 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_888 = _T_63 ? _GEN_849 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_889 = _T_63 ? _GEN_850 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_890 = _T_63 ? _GEN_851 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_891 = _T_63 ? _GEN_852 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_892 = _T_63 ? _GEN_853 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_893 = _T_63 ? _GEN_854 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_894 = _T_63 ? _GEN_855 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_895 = _T_63 ? _GEN_856 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_896 = _T_63 ? _GEN_857 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_897 = _T_63 ? _GEN_858 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_898 = _T_63 ? _GEN_859 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_899 = _T_63 ? _GEN_860 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_900 = _T_63 ? _GEN_861 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_901 = _T_63 ? _GEN_862 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_902 = _T_63 ? _GEN_863 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_903 = _T_63 ? _GEN_864 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_904 = _T_63 ? _GEN_865 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_905 = _T_63 ? _GEN_866 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_906 = _T_63 ? _GEN_867 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_907 = _T_63 ? _GEN_868 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_908 = _T_63 ? _GEN_869 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_909 = _T_63 ? _GEN_870 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_910 = _T_63 ? _GEN_871 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [31:0] _GEN_911 = _T_63 ? _GEN_872 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [6:0] _funct7_T_1 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_10 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_75 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_9 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_23 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:66]
  wire [31:0] _now_reg_rs2_0 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_24 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:88]
  wire  _next_reg_T_25 = $signed(_T_300) < $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:73]
  wire  _next_reg_T_26 = _T_246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:73]
  wire [31:0] _next_reg_rd_11 = {{31'd0}, _T_246}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_912 = 5'h0 == rd ? _next_reg_rd_11 : _GEN_880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_913 = 5'h1 == rd ? _next_reg_rd_11 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_914 = 5'h2 == rd ? _next_reg_rd_11 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_915 = 5'h3 == rd ? _next_reg_rd_11 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_916 = 5'h4 == rd ? _next_reg_rd_11 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_917 = 5'h5 == rd ? _next_reg_rd_11 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_918 = 5'h6 == rd ? _next_reg_rd_11 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_919 = 5'h7 == rd ? _next_reg_rd_11 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_920 = 5'h8 == rd ? _next_reg_rd_11 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_921 = 5'h9 == rd ? _next_reg_rd_11 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_922 = 5'ha == rd ? _next_reg_rd_11 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_923 = 5'hb == rd ? _next_reg_rd_11 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_924 = 5'hc == rd ? _next_reg_rd_11 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_925 = 5'hd == rd ? _next_reg_rd_11 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_926 = 5'he == rd ? _next_reg_rd_11 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_927 = 5'hf == rd ? _next_reg_rd_11 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_928 = 5'h10 == rd ? _next_reg_rd_11 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_929 = 5'h11 == rd ? _next_reg_rd_11 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_930 = 5'h12 == rd ? _next_reg_rd_11 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_931 = 5'h13 == rd ? _next_reg_rd_11 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_932 = 5'h14 == rd ? _next_reg_rd_11 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_933 = 5'h15 == rd ? _next_reg_rd_11 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_934 = 5'h16 == rd ? _next_reg_rd_11 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_935 = 5'h17 == rd ? _next_reg_rd_11 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_936 = 5'h18 == rd ? _next_reg_rd_11 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_937 = 5'h19 == rd ? _next_reg_rd_11 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_938 = 5'h1a == rd ? _next_reg_rd_11 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_939 = 5'h1b == rd ? _next_reg_rd_11 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_940 = 5'h1c == rd ? _next_reg_rd_11 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_941 = 5'h1d == rd ? _next_reg_rd_11 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_942 = 5'h1e == rd ? _next_reg_rd_11 : _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [31:0] _GEN_943 = 5'h1f == rd ? _next_reg_rd_11 : _GEN_911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [6:0] _GEN_945 = _T_70 ? inst[31:25] : _GEN_874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_948 = _T_70 ? inst[14:12] : _GEN_877; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_950 = _T_70 ? inst[6:0] : _GEN_879; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_951 = _T_70 ? _GEN_912 : _GEN_880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_952 = _T_70 ? _GEN_913 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_953 = _T_70 ? _GEN_914 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_954 = _T_70 ? _GEN_915 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_955 = _T_70 ? _GEN_916 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_956 = _T_70 ? _GEN_917 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_957 = _T_70 ? _GEN_918 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_958 = _T_70 ? _GEN_919 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_959 = _T_70 ? _GEN_920 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_960 = _T_70 ? _GEN_921 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_961 = _T_70 ? _GEN_922 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_962 = _T_70 ? _GEN_923 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_963 = _T_70 ? _GEN_924 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_964 = _T_70 ? _GEN_925 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_965 = _T_70 ? _GEN_926 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_966 = _T_70 ? _GEN_927 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_967 = _T_70 ? _GEN_928 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_968 = _T_70 ? _GEN_929 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_969 = _T_70 ? _GEN_930 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_970 = _T_70 ? _GEN_931 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_971 = _T_70 ? _GEN_932 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_972 = _T_70 ? _GEN_933 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_973 = _T_70 ? _GEN_934 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_974 = _T_70 ? _GEN_935 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_975 = _T_70 ? _GEN_936 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_976 = _T_70 ? _GEN_937 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_977 = _T_70 ? _GEN_938 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_978 = _T_70 ? _GEN_939 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_979 = _T_70 ? _GEN_940 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_980 = _T_70 ? _GEN_941 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_981 = _T_70 ? _GEN_942 : _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [31:0] _GEN_982 = _T_70 ? _GEN_943 : _GEN_911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [6:0] _funct7_T_2 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_11 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_82 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_10 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_1 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_27 = _GEN_31 < _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:66]
  wire  _next_reg_T_28 = _T_273; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:66]
  wire [31:0] _next_reg_rd_12 = {{31'd0}, _T_273}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_983 = 5'h0 == rd ? _next_reg_rd_12 : _GEN_951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_984 = 5'h1 == rd ? _next_reg_rd_12 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_985 = 5'h2 == rd ? _next_reg_rd_12 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_986 = 5'h3 == rd ? _next_reg_rd_12 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_987 = 5'h4 == rd ? _next_reg_rd_12 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_988 = 5'h5 == rd ? _next_reg_rd_12 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_989 = 5'h6 == rd ? _next_reg_rd_12 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_990 = 5'h7 == rd ? _next_reg_rd_12 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_991 = 5'h8 == rd ? _next_reg_rd_12 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_992 = 5'h9 == rd ? _next_reg_rd_12 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_993 = 5'ha == rd ? _next_reg_rd_12 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_994 = 5'hb == rd ? _next_reg_rd_12 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_995 = 5'hc == rd ? _next_reg_rd_12 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_996 = 5'hd == rd ? _next_reg_rd_12 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_997 = 5'he == rd ? _next_reg_rd_12 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_998 = 5'hf == rd ? _next_reg_rd_12 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_999 = 5'h10 == rd ? _next_reg_rd_12 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1000 = 5'h11 == rd ? _next_reg_rd_12 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1001 = 5'h12 == rd ? _next_reg_rd_12 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1002 = 5'h13 == rd ? _next_reg_rd_12 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1003 = 5'h14 == rd ? _next_reg_rd_12 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1004 = 5'h15 == rd ? _next_reg_rd_12 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1005 = 5'h16 == rd ? _next_reg_rd_12 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1006 = 5'h17 == rd ? _next_reg_rd_12 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1007 = 5'h18 == rd ? _next_reg_rd_12 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1008 = 5'h19 == rd ? _next_reg_rd_12 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1009 = 5'h1a == rd ? _next_reg_rd_12 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1010 = 5'h1b == rd ? _next_reg_rd_12 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1011 = 5'h1c == rd ? _next_reg_rd_12 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1012 = 5'h1d == rd ? _next_reg_rd_12 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1013 = 5'h1e == rd ? _next_reg_rd_12 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [31:0] _GEN_1014 = 5'h1f == rd ? _next_reg_rd_12 : _GEN_982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [6:0] _GEN_1016 = _T_77 ? inst[31:25] : _GEN_945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1019 = _T_77 ? inst[14:12] : _GEN_948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1021 = _T_77 ? inst[6:0] : _GEN_950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1022 = _T_77 ? _GEN_983 : _GEN_951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1023 = _T_77 ? _GEN_984 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1024 = _T_77 ? _GEN_985 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1025 = _T_77 ? _GEN_986 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1026 = _T_77 ? _GEN_987 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1027 = _T_77 ? _GEN_988 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1028 = _T_77 ? _GEN_989 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1029 = _T_77 ? _GEN_990 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1030 = _T_77 ? _GEN_991 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1031 = _T_77 ? _GEN_992 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1032 = _T_77 ? _GEN_993 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1033 = _T_77 ? _GEN_994 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1034 = _T_77 ? _GEN_995 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1035 = _T_77 ? _GEN_996 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1036 = _T_77 ? _GEN_997 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1037 = _T_77 ? _GEN_998 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1038 = _T_77 ? _GEN_999 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1039 = _T_77 ? _GEN_1000 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1040 = _T_77 ? _GEN_1001 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1041 = _T_77 ? _GEN_1002 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1042 = _T_77 ? _GEN_1003 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1043 = _T_77 ? _GEN_1004 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1044 = _T_77 ? _GEN_1005 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1045 = _T_77 ? _GEN_1006 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1046 = _T_77 ? _GEN_1007 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1047 = _T_77 ? _GEN_1008 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1048 = _T_77 ? _GEN_1009 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1049 = _T_77 ? _GEN_1010 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1050 = _T_77 ? _GEN_1011 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1051 = _T_77 ? _GEN_1012 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1052 = _T_77 ? _GEN_1013 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [31:0] _GEN_1053 = _T_77 ? _GEN_1014 : _GEN_982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [6:0] _funct7_T_3 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_12 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_89 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_11 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_2 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_29 = _GEN_31 & _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:61]
  wire [31:0] _next_reg_rd_13 = _GEN_31 & _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:61]
  wire [31:0] _GEN_1054 = 5'h0 == rd ? _next_reg_T_29 : _GEN_1022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1055 = 5'h1 == rd ? _next_reg_T_29 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1056 = 5'h2 == rd ? _next_reg_T_29 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1057 = 5'h3 == rd ? _next_reg_T_29 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1058 = 5'h4 == rd ? _next_reg_T_29 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1059 = 5'h5 == rd ? _next_reg_T_29 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1060 = 5'h6 == rd ? _next_reg_T_29 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1061 = 5'h7 == rd ? _next_reg_T_29 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1062 = 5'h8 == rd ? _next_reg_T_29 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1063 = 5'h9 == rd ? _next_reg_T_29 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1064 = 5'ha == rd ? _next_reg_T_29 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1065 = 5'hb == rd ? _next_reg_T_29 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1066 = 5'hc == rd ? _next_reg_T_29 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1067 = 5'hd == rd ? _next_reg_T_29 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1068 = 5'he == rd ? _next_reg_T_29 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1069 = 5'hf == rd ? _next_reg_T_29 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1070 = 5'h10 == rd ? _next_reg_T_29 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1071 = 5'h11 == rd ? _next_reg_T_29 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1072 = 5'h12 == rd ? _next_reg_T_29 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1073 = 5'h13 == rd ? _next_reg_T_29 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1074 = 5'h14 == rd ? _next_reg_T_29 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1075 = 5'h15 == rd ? _next_reg_T_29 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1076 = 5'h16 == rd ? _next_reg_T_29 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1077 = 5'h17 == rd ? _next_reg_T_29 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1078 = 5'h18 == rd ? _next_reg_T_29 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1079 = 5'h19 == rd ? _next_reg_T_29 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1080 = 5'h1a == rd ? _next_reg_T_29 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1081 = 5'h1b == rd ? _next_reg_T_29 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1082 = 5'h1c == rd ? _next_reg_T_29 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1083 = 5'h1d == rd ? _next_reg_T_29 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1084 = 5'h1e == rd ? _next_reg_T_29 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [31:0] _GEN_1085 = 5'h1f == rd ? _next_reg_T_29 : _GEN_1053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [6:0] _GEN_1087 = _T_84 ? inst[31:25] : _GEN_1016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1090 = _T_84 ? inst[14:12] : _GEN_1019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1092 = _T_84 ? inst[6:0] : _GEN_1021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1093 = _T_84 ? _GEN_1054 : _GEN_1022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1094 = _T_84 ? _GEN_1055 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1095 = _T_84 ? _GEN_1056 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1096 = _T_84 ? _GEN_1057 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1097 = _T_84 ? _GEN_1058 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1098 = _T_84 ? _GEN_1059 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1099 = _T_84 ? _GEN_1060 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1100 = _T_84 ? _GEN_1061 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1101 = _T_84 ? _GEN_1062 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1102 = _T_84 ? _GEN_1063 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1103 = _T_84 ? _GEN_1064 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1104 = _T_84 ? _GEN_1065 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1105 = _T_84 ? _GEN_1066 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1106 = _T_84 ? _GEN_1067 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1107 = _T_84 ? _GEN_1068 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1108 = _T_84 ? _GEN_1069 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1109 = _T_84 ? _GEN_1070 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1110 = _T_84 ? _GEN_1071 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1111 = _T_84 ? _GEN_1072 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1112 = _T_84 ? _GEN_1073 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1113 = _T_84 ? _GEN_1074 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1114 = _T_84 ? _GEN_1075 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1115 = _T_84 ? _GEN_1076 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1116 = _T_84 ? _GEN_1077 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1117 = _T_84 ? _GEN_1078 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1118 = _T_84 ? _GEN_1079 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1119 = _T_84 ? _GEN_1080 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1120 = _T_84 ? _GEN_1081 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1121 = _T_84 ? _GEN_1082 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1122 = _T_84 ? _GEN_1083 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1123 = _T_84 ? _GEN_1084 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [31:0] _GEN_1124 = _T_84 ? _GEN_1085 : _GEN_1053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [6:0] _funct7_T_4 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_13 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_96 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_12 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_3 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_30 = _GEN_31 | _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:61]
  wire [31:0] _next_reg_rd_14 = _GEN_31 | _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:61]
  wire [31:0] _GEN_1125 = 5'h0 == rd ? _next_reg_T_30 : _GEN_1093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1126 = 5'h1 == rd ? _next_reg_T_30 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1127 = 5'h2 == rd ? _next_reg_T_30 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1128 = 5'h3 == rd ? _next_reg_T_30 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1129 = 5'h4 == rd ? _next_reg_T_30 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1130 = 5'h5 == rd ? _next_reg_T_30 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1131 = 5'h6 == rd ? _next_reg_T_30 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1132 = 5'h7 == rd ? _next_reg_T_30 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1133 = 5'h8 == rd ? _next_reg_T_30 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1134 = 5'h9 == rd ? _next_reg_T_30 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1135 = 5'ha == rd ? _next_reg_T_30 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1136 = 5'hb == rd ? _next_reg_T_30 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1137 = 5'hc == rd ? _next_reg_T_30 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1138 = 5'hd == rd ? _next_reg_T_30 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1139 = 5'he == rd ? _next_reg_T_30 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1140 = 5'hf == rd ? _next_reg_T_30 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1141 = 5'h10 == rd ? _next_reg_T_30 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1142 = 5'h11 == rd ? _next_reg_T_30 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1143 = 5'h12 == rd ? _next_reg_T_30 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1144 = 5'h13 == rd ? _next_reg_T_30 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1145 = 5'h14 == rd ? _next_reg_T_30 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1146 = 5'h15 == rd ? _next_reg_T_30 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1147 = 5'h16 == rd ? _next_reg_T_30 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1148 = 5'h17 == rd ? _next_reg_T_30 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1149 = 5'h18 == rd ? _next_reg_T_30 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1150 = 5'h19 == rd ? _next_reg_T_30 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1151 = 5'h1a == rd ? _next_reg_T_30 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1152 = 5'h1b == rd ? _next_reg_T_30 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1153 = 5'h1c == rd ? _next_reg_T_30 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1154 = 5'h1d == rd ? _next_reg_T_30 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1155 = 5'h1e == rd ? _next_reg_T_30 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [31:0] _GEN_1156 = 5'h1f == rd ? _next_reg_T_30 : _GEN_1124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [6:0] _GEN_1158 = _T_91 ? inst[31:25] : _GEN_1087; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1161 = _T_91 ? inst[14:12] : _GEN_1090; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1163 = _T_91 ? inst[6:0] : _GEN_1092; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1164 = _T_91 ? _GEN_1125 : _GEN_1093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1165 = _T_91 ? _GEN_1126 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1166 = _T_91 ? _GEN_1127 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1167 = _T_91 ? _GEN_1128 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1168 = _T_91 ? _GEN_1129 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1169 = _T_91 ? _GEN_1130 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1170 = _T_91 ? _GEN_1131 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1171 = _T_91 ? _GEN_1132 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1172 = _T_91 ? _GEN_1133 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1173 = _T_91 ? _GEN_1134 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1174 = _T_91 ? _GEN_1135 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1175 = _T_91 ? _GEN_1136 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1176 = _T_91 ? _GEN_1137 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1177 = _T_91 ? _GEN_1138 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1178 = _T_91 ? _GEN_1139 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1179 = _T_91 ? _GEN_1140 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1180 = _T_91 ? _GEN_1141 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1181 = _T_91 ? _GEN_1142 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1182 = _T_91 ? _GEN_1143 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1183 = _T_91 ? _GEN_1144 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1184 = _T_91 ? _GEN_1145 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1185 = _T_91 ? _GEN_1146 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1186 = _T_91 ? _GEN_1147 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1187 = _T_91 ? _GEN_1148 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1188 = _T_91 ? _GEN_1149 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1189 = _T_91 ? _GEN_1150 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1190 = _T_91 ? _GEN_1151 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1191 = _T_91 ? _GEN_1152 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1192 = _T_91 ? _GEN_1153 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1193 = _T_91 ? _GEN_1154 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1194 = _T_91 ? _GEN_1155 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [31:0] _GEN_1195 = _T_91 ? _GEN_1156 : _GEN_1124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [6:0] _funct7_T_5 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_14 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_103 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_13 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_4 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_31 = _GEN_31 ^ _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:61]
  wire [31:0] _next_reg_rd_15 = _GEN_31 ^ _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:61]
  wire [31:0] _GEN_1196 = 5'h0 == rd ? _next_reg_T_31 : _GEN_1164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1197 = 5'h1 == rd ? _next_reg_T_31 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1198 = 5'h2 == rd ? _next_reg_T_31 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1199 = 5'h3 == rd ? _next_reg_T_31 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1200 = 5'h4 == rd ? _next_reg_T_31 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1201 = 5'h5 == rd ? _next_reg_T_31 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1202 = 5'h6 == rd ? _next_reg_T_31 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1203 = 5'h7 == rd ? _next_reg_T_31 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1204 = 5'h8 == rd ? _next_reg_T_31 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1205 = 5'h9 == rd ? _next_reg_T_31 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1206 = 5'ha == rd ? _next_reg_T_31 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1207 = 5'hb == rd ? _next_reg_T_31 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1208 = 5'hc == rd ? _next_reg_T_31 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1209 = 5'hd == rd ? _next_reg_T_31 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1210 = 5'he == rd ? _next_reg_T_31 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1211 = 5'hf == rd ? _next_reg_T_31 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1212 = 5'h10 == rd ? _next_reg_T_31 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1213 = 5'h11 == rd ? _next_reg_T_31 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1214 = 5'h12 == rd ? _next_reg_T_31 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1215 = 5'h13 == rd ? _next_reg_T_31 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1216 = 5'h14 == rd ? _next_reg_T_31 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1217 = 5'h15 == rd ? _next_reg_T_31 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1218 = 5'h16 == rd ? _next_reg_T_31 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1219 = 5'h17 == rd ? _next_reg_T_31 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1220 = 5'h18 == rd ? _next_reg_T_31 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1221 = 5'h19 == rd ? _next_reg_T_31 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1222 = 5'h1a == rd ? _next_reg_T_31 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1223 = 5'h1b == rd ? _next_reg_T_31 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1224 = 5'h1c == rd ? _next_reg_T_31 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1225 = 5'h1d == rd ? _next_reg_T_31 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1226 = 5'h1e == rd ? _next_reg_T_31 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [31:0] _GEN_1227 = 5'h1f == rd ? _next_reg_T_31 : _GEN_1195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [6:0] _GEN_1229 = _T_98 ? inst[31:25] : _GEN_1158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1232 = _T_98 ? inst[14:12] : _GEN_1161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1234 = _T_98 ? inst[6:0] : _GEN_1163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1235 = _T_98 ? _GEN_1196 : _GEN_1164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1236 = _T_98 ? _GEN_1197 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1237 = _T_98 ? _GEN_1198 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1238 = _T_98 ? _GEN_1199 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1239 = _T_98 ? _GEN_1200 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1240 = _T_98 ? _GEN_1201 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1241 = _T_98 ? _GEN_1202 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1242 = _T_98 ? _GEN_1203 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1243 = _T_98 ? _GEN_1204 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1244 = _T_98 ? _GEN_1205 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1245 = _T_98 ? _GEN_1206 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1246 = _T_98 ? _GEN_1207 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1247 = _T_98 ? _GEN_1208 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1248 = _T_98 ? _GEN_1209 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1249 = _T_98 ? _GEN_1210 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1250 = _T_98 ? _GEN_1211 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1251 = _T_98 ? _GEN_1212 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1252 = _T_98 ? _GEN_1213 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1253 = _T_98 ? _GEN_1214 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1254 = _T_98 ? _GEN_1215 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1255 = _T_98 ? _GEN_1216 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1256 = _T_98 ? _GEN_1217 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1257 = _T_98 ? _GEN_1218 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1258 = _T_98 ? _GEN_1219 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1259 = _T_98 ? _GEN_1220 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1260 = _T_98 ? _GEN_1221 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1261 = _T_98 ? _GEN_1222 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1262 = _T_98 ? _GEN_1223 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1263 = _T_98 ? _GEN_1224 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1264 = _T_98 ? _GEN_1225 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1265 = _T_98 ? _GEN_1226 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [31:0] _GEN_1266 = _T_98 ? _GEN_1227 : _GEN_1195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [6:0] _funct7_T_6 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_15 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_110 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs2_5 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [4:0] _next_reg_T_32 = _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:76]
  wire [31:0] _now_reg_rs1_14 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [62:0] _GEN_3348 = {{31'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [62:0] _next_reg_T_33 = _GEN_3348 << _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [31:0] _next_reg_rd_16 = _next_reg_T_33[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1267 = 5'h0 == rd ? _next_reg_T_33[31:0] : _GEN_1235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1268 = 5'h1 == rd ? _next_reg_T_33[31:0] : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1269 = 5'h2 == rd ? _next_reg_T_33[31:0] : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1270 = 5'h3 == rd ? _next_reg_T_33[31:0] : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1271 = 5'h4 == rd ? _next_reg_T_33[31:0] : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1272 = 5'h5 == rd ? _next_reg_T_33[31:0] : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1273 = 5'h6 == rd ? _next_reg_T_33[31:0] : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1274 = 5'h7 == rd ? _next_reg_T_33[31:0] : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1275 = 5'h8 == rd ? _next_reg_T_33[31:0] : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1276 = 5'h9 == rd ? _next_reg_T_33[31:0] : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1277 = 5'ha == rd ? _next_reg_T_33[31:0] : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1278 = 5'hb == rd ? _next_reg_T_33[31:0] : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1279 = 5'hc == rd ? _next_reg_T_33[31:0] : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1280 = 5'hd == rd ? _next_reg_T_33[31:0] : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1281 = 5'he == rd ? _next_reg_T_33[31:0] : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1282 = 5'hf == rd ? _next_reg_T_33[31:0] : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1283 = 5'h10 == rd ? _next_reg_T_33[31:0] : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1284 = 5'h11 == rd ? _next_reg_T_33[31:0] : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1285 = 5'h12 == rd ? _next_reg_T_33[31:0] : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1286 = 5'h13 == rd ? _next_reg_T_33[31:0] : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1287 = 5'h14 == rd ? _next_reg_T_33[31:0] : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1288 = 5'h15 == rd ? _next_reg_T_33[31:0] : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1289 = 5'h16 == rd ? _next_reg_T_33[31:0] : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1290 = 5'h17 == rd ? _next_reg_T_33[31:0] : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1291 = 5'h18 == rd ? _next_reg_T_33[31:0] : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1292 = 5'h19 == rd ? _next_reg_T_33[31:0] : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1293 = 5'h1a == rd ? _next_reg_T_33[31:0] : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1294 = 5'h1b == rd ? _next_reg_T_33[31:0] : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1295 = 5'h1c == rd ? _next_reg_T_33[31:0] : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1296 = 5'h1d == rd ? _next_reg_T_33[31:0] : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1297 = 5'h1e == rd ? _next_reg_T_33[31:0] : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [31:0] _GEN_1298 = 5'h1f == rd ? _next_reg_T_33[31:0] : _GEN_1266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [6:0] _GEN_1300 = _T_105 ? inst[31:25] : _GEN_1229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1303 = _T_105 ? inst[14:12] : _GEN_1232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1305 = _T_105 ? inst[6:0] : _GEN_1234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1306 = _T_105 ? _GEN_1267 : _GEN_1235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1307 = _T_105 ? _GEN_1268 : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1308 = _T_105 ? _GEN_1269 : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1309 = _T_105 ? _GEN_1270 : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1310 = _T_105 ? _GEN_1271 : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1311 = _T_105 ? _GEN_1272 : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1312 = _T_105 ? _GEN_1273 : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1313 = _T_105 ? _GEN_1274 : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1314 = _T_105 ? _GEN_1275 : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1315 = _T_105 ? _GEN_1276 : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1316 = _T_105 ? _GEN_1277 : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1317 = _T_105 ? _GEN_1278 : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1318 = _T_105 ? _GEN_1279 : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1319 = _T_105 ? _GEN_1280 : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1320 = _T_105 ? _GEN_1281 : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1321 = _T_105 ? _GEN_1282 : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1322 = _T_105 ? _GEN_1283 : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1323 = _T_105 ? _GEN_1284 : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1324 = _T_105 ? _GEN_1285 : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1325 = _T_105 ? _GEN_1286 : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1326 = _T_105 ? _GEN_1287 : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1327 = _T_105 ? _GEN_1288 : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1328 = _T_105 ? _GEN_1289 : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1329 = _T_105 ? _GEN_1290 : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1330 = _T_105 ? _GEN_1291 : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1331 = _T_105 ? _GEN_1292 : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1332 = _T_105 ? _GEN_1293 : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1333 = _T_105 ? _GEN_1294 : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1334 = _T_105 ? _GEN_1295 : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1335 = _T_105 ? _GEN_1296 : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1336 = _T_105 ? _GEN_1297 : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [31:0] _GEN_1337 = _T_105 ? _GEN_1298 : _GEN_1266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [6:0] _funct7_T_7 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_16 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_117 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs2_6 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [4:0] _next_reg_T_34 = _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:76]
  wire [31:0] _now_reg_rs1_15 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_35 = _GEN_31 >> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:61]
  wire [31:0] _next_reg_rd_17 = _GEN_31 >> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:61]
  wire [31:0] _GEN_1338 = 5'h0 == rd ? _next_reg_T_35 : _GEN_1306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1339 = 5'h1 == rd ? _next_reg_T_35 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1340 = 5'h2 == rd ? _next_reg_T_35 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1341 = 5'h3 == rd ? _next_reg_T_35 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1342 = 5'h4 == rd ? _next_reg_T_35 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1343 = 5'h5 == rd ? _next_reg_T_35 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1344 = 5'h6 == rd ? _next_reg_T_35 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1345 = 5'h7 == rd ? _next_reg_T_35 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1346 = 5'h8 == rd ? _next_reg_T_35 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1347 = 5'h9 == rd ? _next_reg_T_35 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1348 = 5'ha == rd ? _next_reg_T_35 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1349 = 5'hb == rd ? _next_reg_T_35 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1350 = 5'hc == rd ? _next_reg_T_35 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1351 = 5'hd == rd ? _next_reg_T_35 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1352 = 5'he == rd ? _next_reg_T_35 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1353 = 5'hf == rd ? _next_reg_T_35 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1354 = 5'h10 == rd ? _next_reg_T_35 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1355 = 5'h11 == rd ? _next_reg_T_35 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1356 = 5'h12 == rd ? _next_reg_T_35 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1357 = 5'h13 == rd ? _next_reg_T_35 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1358 = 5'h14 == rd ? _next_reg_T_35 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1359 = 5'h15 == rd ? _next_reg_T_35 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1360 = 5'h16 == rd ? _next_reg_T_35 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1361 = 5'h17 == rd ? _next_reg_T_35 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1362 = 5'h18 == rd ? _next_reg_T_35 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1363 = 5'h19 == rd ? _next_reg_T_35 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1364 = 5'h1a == rd ? _next_reg_T_35 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1365 = 5'h1b == rd ? _next_reg_T_35 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1366 = 5'h1c == rd ? _next_reg_T_35 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1367 = 5'h1d == rd ? _next_reg_T_35 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1368 = 5'h1e == rd ? _next_reg_T_35 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [31:0] _GEN_1369 = 5'h1f == rd ? _next_reg_T_35 : _GEN_1337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [6:0] _GEN_1371 = _T_112 ? inst[31:25] : _GEN_1300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1374 = _T_112 ? inst[14:12] : _GEN_1303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1376 = _T_112 ? inst[6:0] : _GEN_1305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1377 = _T_112 ? _GEN_1338 : _GEN_1306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1378 = _T_112 ? _GEN_1339 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1379 = _T_112 ? _GEN_1340 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1380 = _T_112 ? _GEN_1341 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1381 = _T_112 ? _GEN_1342 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1382 = _T_112 ? _GEN_1343 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1383 = _T_112 ? _GEN_1344 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1384 = _T_112 ? _GEN_1345 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1385 = _T_112 ? _GEN_1346 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1386 = _T_112 ? _GEN_1347 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1387 = _T_112 ? _GEN_1348 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1388 = _T_112 ? _GEN_1349 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1389 = _T_112 ? _GEN_1350 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1390 = _T_112 ? _GEN_1351 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1391 = _T_112 ? _GEN_1352 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1392 = _T_112 ? _GEN_1353 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1393 = _T_112 ? _GEN_1354 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1394 = _T_112 ? _GEN_1355 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1395 = _T_112 ? _GEN_1356 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1396 = _T_112 ? _GEN_1357 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1397 = _T_112 ? _GEN_1358 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1398 = _T_112 ? _GEN_1359 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1399 = _T_112 ? _GEN_1360 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1400 = _T_112 ? _GEN_1361 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1401 = _T_112 ? _GEN_1362 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1402 = _T_112 ? _GEN_1363 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1403 = _T_112 ? _GEN_1364 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1404 = _T_112 ? _GEN_1365 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1405 = _T_112 ? _GEN_1366 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1406 = _T_112 ? _GEN_1367 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1407 = _T_112 ? _GEN_1368 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [31:0] _GEN_1408 = _T_112 ? _GEN_1369 : _GEN_1337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [6:0] _funct7_T_8 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_17 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_124 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_16 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_7 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_36 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [31:0] _next_reg_T_37 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [31:0] _next_reg_rd_18 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [31:0] _GEN_1409 = 5'h0 == rd ? _next_reg_T_37 : _GEN_1377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1410 = 5'h1 == rd ? _next_reg_T_37 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1411 = 5'h2 == rd ? _next_reg_T_37 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1412 = 5'h3 == rd ? _next_reg_T_37 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1413 = 5'h4 == rd ? _next_reg_T_37 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1414 = 5'h5 == rd ? _next_reg_T_37 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1415 = 5'h6 == rd ? _next_reg_T_37 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1416 = 5'h7 == rd ? _next_reg_T_37 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1417 = 5'h8 == rd ? _next_reg_T_37 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1418 = 5'h9 == rd ? _next_reg_T_37 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1419 = 5'ha == rd ? _next_reg_T_37 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1420 = 5'hb == rd ? _next_reg_T_37 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1421 = 5'hc == rd ? _next_reg_T_37 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1422 = 5'hd == rd ? _next_reg_T_37 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1423 = 5'he == rd ? _next_reg_T_37 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1424 = 5'hf == rd ? _next_reg_T_37 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1425 = 5'h10 == rd ? _next_reg_T_37 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1426 = 5'h11 == rd ? _next_reg_T_37 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1427 = 5'h12 == rd ? _next_reg_T_37 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1428 = 5'h13 == rd ? _next_reg_T_37 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1429 = 5'h14 == rd ? _next_reg_T_37 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1430 = 5'h15 == rd ? _next_reg_T_37 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1431 = 5'h16 == rd ? _next_reg_T_37 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1432 = 5'h17 == rd ? _next_reg_T_37 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1433 = 5'h18 == rd ? _next_reg_T_37 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1434 = 5'h19 == rd ? _next_reg_T_37 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1435 = 5'h1a == rd ? _next_reg_T_37 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1436 = 5'h1b == rd ? _next_reg_T_37 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1437 = 5'h1c == rd ? _next_reg_T_37 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1438 = 5'h1d == rd ? _next_reg_T_37 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1439 = 5'h1e == rd ? _next_reg_T_37 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [31:0] _GEN_1440 = 5'h1f == rd ? _next_reg_T_37 : _GEN_1408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [6:0] _GEN_1442 = _T_119 ? inst[31:25] : _GEN_1371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1445 = _T_119 ? inst[14:12] : _GEN_1374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1447 = _T_119 ? inst[6:0] : _GEN_1376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1448 = _T_119 ? _GEN_1409 : _GEN_1377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1449 = _T_119 ? _GEN_1410 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1450 = _T_119 ? _GEN_1411 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1451 = _T_119 ? _GEN_1412 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1452 = _T_119 ? _GEN_1413 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1453 = _T_119 ? _GEN_1414 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1454 = _T_119 ? _GEN_1415 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1455 = _T_119 ? _GEN_1416 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1456 = _T_119 ? _GEN_1417 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1457 = _T_119 ? _GEN_1418 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1458 = _T_119 ? _GEN_1419 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1459 = _T_119 ? _GEN_1420 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1460 = _T_119 ? _GEN_1421 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1461 = _T_119 ? _GEN_1422 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1462 = _T_119 ? _GEN_1423 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1463 = _T_119 ? _GEN_1424 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1464 = _T_119 ? _GEN_1425 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1465 = _T_119 ? _GEN_1426 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1466 = _T_119 ? _GEN_1427 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1467 = _T_119 ? _GEN_1428 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1468 = _T_119 ? _GEN_1429 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1469 = _T_119 ? _GEN_1430 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1470 = _T_119 ? _GEN_1431 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1471 = _T_119 ? _GEN_1432 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1472 = _T_119 ? _GEN_1433 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1473 = _T_119 ? _GEN_1434 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1474 = _T_119 ? _GEN_1435 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1475 = _T_119 ? _GEN_1436 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1476 = _T_119 ? _GEN_1437 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1477 = _T_119 ? _GEN_1438 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1478 = _T_119 ? _GEN_1439 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [31:0] _GEN_1479 = _T_119 ? _GEN_1440 : _GEN_1408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [6:0] _funct7_T_9 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_18 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_131 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_17 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_38 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:62]
  wire [31:0] _now_reg_rs2_8 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [4:0] _next_reg_T_39 = _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:84]
  wire [31:0] _next_reg_T_40 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:69]
  wire [31:0] _next_reg_T_41 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:92]
  wire [31:0] _next_reg_rd_19 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:92]
  wire [31:0] _GEN_1480 = 5'h0 == rd ? _next_reg_T_41 : _GEN_1448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1481 = 5'h1 == rd ? _next_reg_T_41 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1482 = 5'h2 == rd ? _next_reg_T_41 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1483 = 5'h3 == rd ? _next_reg_T_41 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1484 = 5'h4 == rd ? _next_reg_T_41 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1485 = 5'h5 == rd ? _next_reg_T_41 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1486 = 5'h6 == rd ? _next_reg_T_41 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1487 = 5'h7 == rd ? _next_reg_T_41 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1488 = 5'h8 == rd ? _next_reg_T_41 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1489 = 5'h9 == rd ? _next_reg_T_41 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1490 = 5'ha == rd ? _next_reg_T_41 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1491 = 5'hb == rd ? _next_reg_T_41 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1492 = 5'hc == rd ? _next_reg_T_41 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1493 = 5'hd == rd ? _next_reg_T_41 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1494 = 5'he == rd ? _next_reg_T_41 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1495 = 5'hf == rd ? _next_reg_T_41 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1496 = 5'h10 == rd ? _next_reg_T_41 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1497 = 5'h11 == rd ? _next_reg_T_41 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1498 = 5'h12 == rd ? _next_reg_T_41 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1499 = 5'h13 == rd ? _next_reg_T_41 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1500 = 5'h14 == rd ? _next_reg_T_41 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1501 = 5'h15 == rd ? _next_reg_T_41 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1502 = 5'h16 == rd ? _next_reg_T_41 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1503 = 5'h17 == rd ? _next_reg_T_41 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1504 = 5'h18 == rd ? _next_reg_T_41 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1505 = 5'h19 == rd ? _next_reg_T_41 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1506 = 5'h1a == rd ? _next_reg_T_41 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1507 = 5'h1b == rd ? _next_reg_T_41 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1508 = 5'h1c == rd ? _next_reg_T_41 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1509 = 5'h1d == rd ? _next_reg_T_41 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1510 = 5'h1e == rd ? _next_reg_T_41 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [31:0] _GEN_1511 = 5'h1f == rd ? _next_reg_T_41 : _GEN_1479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [6:0] _GEN_1513 = _T_126 ? inst[31:25] : _GEN_1442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_1516 = _T_126 ? inst[14:12] : _GEN_1445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1518 = _T_126 ? inst[6:0] : _GEN_1447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_1519 = _T_126 ? _GEN_1480 : _GEN_1448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1520 = _T_126 ? _GEN_1481 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1521 = _T_126 ? _GEN_1482 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1522 = _T_126 ? _GEN_1483 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1523 = _T_126 ? _GEN_1484 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1524 = _T_126 ? _GEN_1485 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1525 = _T_126 ? _GEN_1486 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1526 = _T_126 ? _GEN_1487 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1527 = _T_126 ? _GEN_1488 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1528 = _T_126 ? _GEN_1489 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1529 = _T_126 ? _GEN_1490 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1530 = _T_126 ? _GEN_1491 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1531 = _T_126 ? _GEN_1492 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1532 = _T_126 ? _GEN_1493 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1533 = _T_126 ? _GEN_1494 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1534 = _T_126 ? _GEN_1495 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1535 = _T_126 ? _GEN_1496 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1536 = _T_126 ? _GEN_1497 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1537 = _T_126 ? _GEN_1498 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1538 = _T_126 ? _GEN_1499 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1539 = _T_126 ? _GEN_1500 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1540 = _T_126 ? _GEN_1501 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1541 = _T_126 ? _GEN_1502 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1542 = _T_126 ? _GEN_1503 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1543 = _T_126 ? _GEN_1504 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1544 = _T_126 ? _GEN_1505 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1545 = _T_126 ? _GEN_1506 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1546 = _T_126 ? _GEN_1507 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1547 = _T_126 ? _GEN_1508 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1548 = _T_126 ? _GEN_1509 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1549 = _T_126 ? _GEN_1510 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [31:0] _GEN_1550 = _T_126 ? _GEN_1511 : _GEN_1479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [6:0] _T_138 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 191:37]
  wire [31:0] _next_pc_T_1 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 191:37]
  wire [32:0] _next_reg_T_42 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [31:0] _next_reg_T_43 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [31:0] _next_reg_rd_20 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [31:0] _GEN_1551 = 5'h0 == rd ? _next_reg_T_43 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1552 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1553 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1554 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1555 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1556 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1557 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1558 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1559 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1560 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1561 = 5'ha == rd ? _next_reg_T_43 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1562 = 5'hb == rd ? _next_reg_T_43 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1563 = 5'hc == rd ? _next_reg_T_43 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1564 = 5'hd == rd ? _next_reg_T_43 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1565 = 5'he == rd ? _next_reg_T_43 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1566 = 5'hf == rd ? _next_reg_T_43 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1567 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1568 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1569 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1570 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1571 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1572 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1573 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1574 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1575 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1576 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1577 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1578 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1579 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1580 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1581 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [31:0] _GEN_1582 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [32:0] _next_csr_mtval_T = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 194:34]
  wire [31:0] _next_csr_mtval_T_1 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 194:34]
  wire  _GEN_1583 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [31:0] _GEN_1584 = _T_346 ? _T_334 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 191:27]
  wire [31:0] _GEN_1585 = _T_346 ? _GEN_1551 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1586 = _T_346 ? _GEN_1552 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1587 = _T_346 ? _GEN_1553 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1588 = _T_346 ? _GEN_1554 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1589 = _T_346 ? _GEN_1555 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1590 = _T_346 ? _GEN_1556 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1591 = _T_346 ? _GEN_1557 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1592 = _T_346 ? _GEN_1558 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1593 = _T_346 ? _GEN_1559 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1594 = _T_346 ? _GEN_1560 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1595 = _T_346 ? _GEN_1561 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1596 = _T_346 ? _GEN_1562 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1597 = _T_346 ? _GEN_1563 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1598 = _T_346 ? _GEN_1564 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1599 = _T_346 ? _GEN_1565 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1600 = _T_346 ? _GEN_1566 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1601 = _T_346 ? _GEN_1567 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1602 = _T_346 ? _GEN_1568 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1603 = _T_346 ? _GEN_1569 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1604 = _T_346 ? _GEN_1570 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1605 = _T_346 ? _GEN_1571 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1606 = _T_346 ? _GEN_1572 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1607 = _T_346 ? _GEN_1573 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1608 = _T_346 ? _GEN_1574 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1609 = _T_346 ? _GEN_1575 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1610 = _T_346 ? _GEN_1576 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1611 = _T_346 ? _GEN_1577 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1612 = _T_346 ? _GEN_1578 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1613 = _T_346 ? _GEN_1579 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1614 = _T_346 ? _GEN_1580 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1615 = _T_346 ? _GEN_1581 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] _GEN_1616 = _T_346 ? _GEN_1582 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [31:0] now_csr_mtval = io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_1617 = _T_346 ? io_now_csr_mtval : _T_334; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 194:24]
  wire  _GEN_1619 = _T_346 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36 145:33]
  wire [6:0] _GEN_1626 = _T_133 ? inst[6:0] : _GEN_1518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1628 = _T_133 & _T_346; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 113:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1629 = _T_133 ? _GEN_1584 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1630 = _T_133 ? _GEN_1585 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1631 = _T_133 ? _GEN_1586 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1632 = _T_133 ? _GEN_1587 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1633 = _T_133 ? _GEN_1588 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1634 = _T_133 ? _GEN_1589 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1635 = _T_133 ? _GEN_1590 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1636 = _T_133 ? _GEN_1591 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1637 = _T_133 ? _GEN_1592 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1638 = _T_133 ? _GEN_1593 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1639 = _T_133 ? _GEN_1594 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1640 = _T_133 ? _GEN_1595 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1641 = _T_133 ? _GEN_1596 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1642 = _T_133 ? _GEN_1597 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1643 = _T_133 ? _GEN_1598 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1644 = _T_133 ? _GEN_1599 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1645 = _T_133 ? _GEN_1600 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1646 = _T_133 ? _GEN_1601 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1647 = _T_133 ? _GEN_1602 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1648 = _T_133 ? _GEN_1603 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1649 = _T_133 ? _GEN_1604 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1650 = _T_133 ? _GEN_1605 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1651 = _T_133 ? _GEN_1606 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1652 = _T_133 ? _GEN_1607 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1653 = _T_133 ? _GEN_1608 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1654 = _T_133 ? _GEN_1609 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1655 = _T_133 ? _GEN_1610 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1656 = _T_133 ? _GEN_1611 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1657 = _T_133 ? _GEN_1612 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1658 = _T_133 ? _GEN_1613 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1659 = _T_133 ? _GEN_1614 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1660 = _T_133 ? _GEN_1615 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1661 = _T_133 ? _GEN_1616 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [31:0] _GEN_1662 = _T_133 ? _GEN_1617 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire  _GEN_1664 = _T_133 & _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [2:0] _funct3_T_19 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_161 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_19 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_pc_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:48]
  wire [31:0] _next_pc_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:48]
  wire [30:0] _next_pc_T_4 = _T_433[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:54]
  wire [31:0] _next_pc_T_5 = {_T_433[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 203:33]
  wire [32:0] _next_reg_T_44 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:37]
  wire [31:0] _next_reg_T_45 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:37]
  wire [31:0] _next_reg_rd_21 = _next_reg_T_43; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:37]
  wire [31:0] _GEN_1665 = 5'h0 == rd ? _next_reg_T_43 : _GEN_1630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1666 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1667 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1668 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1669 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1670 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1671 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1672 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1673 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1674 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1675 = 5'ha == rd ? _next_reg_T_43 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1676 = 5'hb == rd ? _next_reg_T_43 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1677 = 5'hc == rd ? _next_reg_T_43 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1678 = 5'hd == rd ? _next_reg_T_43 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1679 = 5'he == rd ? _next_reg_T_43 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1680 = 5'hf == rd ? _next_reg_T_43 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1681 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1682 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1683 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1684 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1685 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1686 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1687 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1688 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1689 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1690 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1691 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1692 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1693 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1694 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1695 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _GEN_1696 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [31:0] _now_reg_rs1_20 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_csr_mtval_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:45]
  wire [31:0] _next_csr_mtval_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:45]
  wire [30:0] _next_csr_mtval_T_4 = _T_433[31:1]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:51]
  wire [31:0] _next_csr_mtval_T_5 = {_T_433[31:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 206:30]
  wire  _GEN_1697 = _T_180 | _GEN_1628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 202:27]
  wire [31:0] _GEN_1698 = _T_180 ? _T_168 : _GEN_1629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 203:27]
  wire [31:0] _GEN_1699 = _T_180 ? _GEN_1665 : _GEN_1630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1700 = _T_180 ? _GEN_1666 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1701 = _T_180 ? _GEN_1667 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1702 = _T_180 ? _GEN_1668 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1703 = _T_180 ? _GEN_1669 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1704 = _T_180 ? _GEN_1670 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1705 = _T_180 ? _GEN_1671 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1706 = _T_180 ? _GEN_1672 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1707 = _T_180 ? _GEN_1673 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1708 = _T_180 ? _GEN_1674 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1709 = _T_180 ? _GEN_1675 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1710 = _T_180 ? _GEN_1676 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1711 = _T_180 ? _GEN_1677 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1712 = _T_180 ? _GEN_1678 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1713 = _T_180 ? _GEN_1679 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1714 = _T_180 ? _GEN_1680 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1715 = _T_180 ? _GEN_1681 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1716 = _T_180 ? _GEN_1682 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1717 = _T_180 ? _GEN_1683 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1718 = _T_180 ? _GEN_1684 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1719 = _T_180 ? _GEN_1685 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1720 = _T_180 ? _GEN_1686 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1721 = _T_180 ? _GEN_1687 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1722 = _T_180 ? _GEN_1688 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1723 = _T_180 ? _GEN_1689 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1724 = _T_180 ? _GEN_1690 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1725 = _T_180 ? _GEN_1691 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1726 = _T_180 ? _GEN_1692 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1727 = _T_180 ? _GEN_1693 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1728 = _T_180 ? _GEN_1694 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1729 = _T_180 ? _GEN_1695 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1730 = _T_180 ? _GEN_1696 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [31:0] _GEN_1731 = _T_180 ? _GEN_1662 : _T_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 206:24]
  wire  _GEN_1733 = _T_180 ? _GEN_1663 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_1737 = _T_157 ? inst[14:12] : _GEN_1516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1739 = _T_157 ? inst[6:0] : _GEN_1626; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1741 = _T_157 ? _GEN_1697 : _GEN_1628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1742 = _T_157 ? _GEN_1698 : _GEN_1629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1743 = _T_157 ? _GEN_1699 : _GEN_1630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1744 = _T_157 ? _GEN_1700 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1745 = _T_157 ? _GEN_1701 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1746 = _T_157 ? _GEN_1702 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1747 = _T_157 ? _GEN_1703 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1748 = _T_157 ? _GEN_1704 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1749 = _T_157 ? _GEN_1705 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1750 = _T_157 ? _GEN_1706 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1751 = _T_157 ? _GEN_1707 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1752 = _T_157 ? _GEN_1708 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1753 = _T_157 ? _GEN_1709 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1754 = _T_157 ? _GEN_1710 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1755 = _T_157 ? _GEN_1711 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1756 = _T_157 ? _GEN_1712 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1757 = _T_157 ? _GEN_1713 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1758 = _T_157 ? _GEN_1714 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1759 = _T_157 ? _GEN_1715 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1760 = _T_157 ? _GEN_1716 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1761 = _T_157 ? _GEN_1717 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1762 = _T_157 ? _GEN_1718 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1763 = _T_157 ? _GEN_1719 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1764 = _T_157 ? _GEN_1720 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1765 = _T_157 ? _GEN_1721 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1766 = _T_157 ? _GEN_1722 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1767 = _T_157 ? _GEN_1723 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1768 = _T_157 ? _GEN_1724 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1769 = _T_157 ? _GEN_1725 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1770 = _T_157 ? _GEN_1726 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1771 = _T_157 ? _GEN_1727 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1772 = _T_157 ? _GEN_1728 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1773 = _T_157 ? _GEN_1729 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1774 = _T_157 ? _GEN_1730 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [31:0] _GEN_1775 = _T_157 ? _GEN_1731 : _GEN_1662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1777 = _T_157 ? _GEN_1732 : _GEN_1663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [2:0] _funct3_T_20 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_189 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_6 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 217:39]
  wire [31:0] _next_pc_T_7 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 217:39]
  wire [32:0] _next_csr_mtval_T_6 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 219:36]
  wire [31:0] _next_csr_mtval_T_7 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 219:36]
  wire  _GEN_1778 = _T_346 | _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 216:29]
  wire [31:0] _GEN_1779 = _T_346 ? _T_334 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 217:29]
  wire [31:0] _GEN_1780 = _T_346 ? _GEN_1775 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 219:26]
  wire  _GEN_1782 = _T_346 ? _GEN_1776 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1783 = _GEN_31 == _GEN_840 ? _GEN_1778 : _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [31:0] _GEN_1784 = _GEN_31 == _GEN_840 ? _GEN_1779 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [31:0] _GEN_1785 = _GEN_31 == _GEN_840 ? _GEN_1780 : _GEN_1775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1787 = _GEN_31 == _GEN_840 ? _GEN_1781 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [2:0] _GEN_1793 = _T_182 ? inst[14:12] : _GEN_1737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1796 = _T_182 ? inst[6:0] : _GEN_1739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1798 = _T_182 ? _GEN_1783 : _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [31:0] _GEN_1799 = _T_182 ? _GEN_1784 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [31:0] _GEN_1800 = _T_182 ? _GEN_1785 : _GEN_1775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1802 = _T_182 ? _GEN_1786 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [2:0] _funct3_T_21 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_216 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_8 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 229:39]
  wire [31:0] _next_pc_T_9 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 229:39]
  wire [32:0] _next_csr_mtval_T_8 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 231:36]
  wire [31:0] _next_csr_mtval_T_9 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 231:36]
  wire  _GEN_1803 = _T_346 | _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 228:29]
  wire [31:0] _GEN_1804 = _T_346 ? _T_334 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 229:29]
  wire [31:0] _GEN_1805 = _T_346 ? _GEN_1800 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 231:26]
  wire  _GEN_1807 = _T_346 ? _GEN_1801 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1808 = _GEN_31 != _GEN_840 ? _GEN_1803 : _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [31:0] _GEN_1809 = _GEN_31 != _GEN_840 ? _GEN_1804 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [31:0] _GEN_1810 = _GEN_31 != _GEN_840 ? _GEN_1805 : _GEN_1800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1812 = _GEN_31 != _GEN_840 ? _GEN_1806 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [2:0] _GEN_1818 = _T_209 ? inst[14:12] : _GEN_1793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1821 = _T_209 ? inst[6:0] : _GEN_1796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1823 = _T_209 ? _GEN_1808 : _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [31:0] _GEN_1824 = _T_209 ? _GEN_1809 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [31:0] _GEN_1825 = _T_209 ? _GEN_1810 : _GEN_1800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1827 = _T_209 ? _GEN_1811 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [2:0] _funct3_T_22 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_243 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_10 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 242:39]
  wire [31:0] _next_pc_T_11 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 242:39]
  wire [32:0] _next_csr_mtval_T_10 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 244:36]
  wire [31:0] _next_csr_mtval_T_11 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 244:36]
  wire  _GEN_1828 = _T_346 | _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 241:29]
  wire [31:0] _GEN_1829 = _T_346 ? _T_334 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 242:29]
  wire [31:0] _GEN_1830 = _T_346 ? _GEN_1825 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 244:26]
  wire  _GEN_1832 = _T_346 ? _GEN_1826 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1833 = $signed(_T_300) < $signed(_T_301) ? _GEN_1828 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [31:0] _GEN_1834 = $signed(_T_300) < $signed(_T_301) ? _GEN_1829 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [31:0] _GEN_1835 = $signed(_T_300) < $signed(_T_301) ? _GEN_1830 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1837 = $signed(_T_300) < $signed(_T_301) ? _GEN_1831 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [2:0] _GEN_1843 = _T_236 ? inst[14:12] : _GEN_1818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1846 = _T_236 ? inst[6:0] : _GEN_1821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1848 = _T_236 ? _GEN_1833 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [31:0] _GEN_1849 = _T_236 ? _GEN_1834 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [31:0] _GEN_1850 = _T_236 ? _GEN_1835 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1852 = _T_236 ? _GEN_1836 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [2:0] _funct3_T_23 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_272 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_12 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 254:39]
  wire [31:0] _next_pc_T_13 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 254:39]
  wire [32:0] _next_csr_mtval_T_12 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 256:36]
  wire [31:0] _next_csr_mtval_T_13 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 256:36]
  wire  _GEN_1853 = _T_346 | _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 253:29]
  wire [31:0] _GEN_1854 = _T_346 ? _T_334 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 254:29]
  wire [31:0] _GEN_1855 = _T_346 ? _GEN_1850 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 256:26]
  wire  _GEN_1857 = _T_346 ? _GEN_1851 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1858 = _GEN_31 < _GEN_840 ? _GEN_1853 : _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [31:0] _GEN_1859 = _GEN_31 < _GEN_840 ? _GEN_1854 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [31:0] _GEN_1860 = _GEN_31 < _GEN_840 ? _GEN_1855 : _GEN_1850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1862 = _GEN_31 < _GEN_840 ? _GEN_1856 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [2:0] _GEN_1868 = _T_265 ? inst[14:12] : _GEN_1843; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1871 = _T_265 ? inst[6:0] : _GEN_1846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1873 = _T_265 ? _GEN_1858 : _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [31:0] _GEN_1874 = _T_265 ? _GEN_1859 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [31:0] _GEN_1875 = _T_265 ? _GEN_1860 : _GEN_1850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1877 = _T_265 ? _GEN_1861 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [2:0] _funct3_T_24 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_299 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_14 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 267:39]
  wire [31:0] _next_pc_T_15 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 267:39]
  wire [32:0] _next_csr_mtval_T_14 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 269:36]
  wire [31:0] _next_csr_mtval_T_15 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 269:36]
  wire  _GEN_1878 = _T_346 | _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 266:29]
  wire [31:0] _GEN_1879 = _T_346 ? _T_334 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 267:29]
  wire [31:0] _GEN_1880 = _T_346 ? _GEN_1875 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 269:26]
  wire  _GEN_1882 = _T_346 ? _GEN_1876 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1883 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1878 : _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [31:0] _GEN_1884 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1879 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [31:0] _GEN_1885 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1880 : _GEN_1875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1887 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1881 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [2:0] _GEN_1893 = _T_292 ? inst[14:12] : _GEN_1868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1896 = _T_292 ? inst[6:0] : _GEN_1871; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1898 = _T_292 ? _GEN_1883 : _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [31:0] _GEN_1899 = _T_292 ? _GEN_1884 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [31:0] _GEN_1900 = _T_292 ? _GEN_1885 : _GEN_1875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1902 = _T_292 ? _GEN_1886 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [2:0] _funct3_T_25 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_328 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [32:0] _next_pc_T_16 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 279:39]
  wire [31:0] _next_pc_T_17 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 279:39]
  wire [32:0] _next_csr_mtval_T_16 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 281:36]
  wire [31:0] _next_csr_mtval_T_17 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 281:36]
  wire  _GEN_1903 = _T_346 | _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 278:29]
  wire [31:0] _GEN_1904 = _T_346 ? _T_334 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 279:29]
  wire [31:0] _GEN_1905 = _T_346 ? _GEN_1900 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 281:26]
  wire  _GEN_1907 = _T_346 ? _GEN_1901 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1908 = _GEN_31 >= _GEN_840 ? _GEN_1903 : _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [31:0] _GEN_1909 = _GEN_31 >= _GEN_840 ? _GEN_1904 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [31:0] _GEN_1910 = _GEN_31 >= _GEN_840 ? _GEN_1905 : _GEN_1900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1912 = _GEN_31 >= _GEN_840 ? _GEN_1906 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [2:0] _GEN_1918 = _T_321 ? inst[14:12] : _GEN_1893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_1921 = _T_321 ? inst[6:0] : _GEN_1896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_1923 = _T_321 ? _GEN_1908 : _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [31:0] _GEN_1924 = _T_321 ? _GEN_1909 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [31:0] _GEN_1925 = _T_321 ? _GEN_1910 : _GEN_1900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  _GEN_1927 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [2:0] _funct3_T_26 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_352 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_28 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_46 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:54]
  wire [31:0] _next_reg_T_47 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:54]
  wire [1:0] _next_reg_rOff_T = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_1 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_2 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_3 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_4 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_5 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_6 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 164:10 21:22]
  wire [31:0] _next_reg_T_48 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_3340 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_49 = _GEN_3340 & 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [7:0] _next_reg_T_50 = _next_reg_T_49[7:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:65]
  wire  next_reg_signBit = _next_reg_T_49[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _next_reg_T_51 = next_reg_signBit; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [23:0] _next_reg_T_52 = next_reg_signBit ? 24'hffffff : 24'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _next_reg_T_53 = {_next_reg_T_52,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _next_reg_rd_22 = {_next_reg_T_52,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_1928 = 5'h0 == rd ? _next_reg_T_53 : _GEN_1743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1929 = 5'h1 == rd ? _next_reg_T_53 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1930 = 5'h2 == rd ? _next_reg_T_53 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1931 = 5'h3 == rd ? _next_reg_T_53 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1932 = 5'h4 == rd ? _next_reg_T_53 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1933 = 5'h5 == rd ? _next_reg_T_53 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1934 = 5'h6 == rd ? _next_reg_T_53 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1935 = 5'h7 == rd ? _next_reg_T_53 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1936 = 5'h8 == rd ? _next_reg_T_53 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1937 = 5'h9 == rd ? _next_reg_T_53 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1938 = 5'ha == rd ? _next_reg_T_53 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1939 = 5'hb == rd ? _next_reg_T_53 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1940 = 5'hc == rd ? _next_reg_T_53 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1941 = 5'hd == rd ? _next_reg_T_53 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1942 = 5'he == rd ? _next_reg_T_53 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1943 = 5'hf == rd ? _next_reg_T_53 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1944 = 5'h10 == rd ? _next_reg_T_53 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1945 = 5'h11 == rd ? _next_reg_T_53 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1946 = 5'h12 == rd ? _next_reg_T_53 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1947 = 5'h13 == rd ? _next_reg_T_53 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1948 = 5'h14 == rd ? _next_reg_T_53 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1949 = 5'h15 == rd ? _next_reg_T_53 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1950 = 5'h16 == rd ? _next_reg_T_53 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1951 = 5'h17 == rd ? _next_reg_T_53 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1952 = 5'h18 == rd ? _next_reg_T_53 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1953 = 5'h19 == rd ? _next_reg_T_53 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1954 = 5'h1a == rd ? _next_reg_T_53 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1955 = 5'h1b == rd ? _next_reg_T_53 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1956 = 5'h1c == rd ? _next_reg_T_53 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1957 = 5'h1d == rd ? _next_reg_T_53 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1958 = 5'h1e == rd ? _next_reg_T_53 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1959 = 5'h1f == rd ? _next_reg_T_53 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _now_reg_rs1_29 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 294:39]
  wire [31:0] _mem_read_addr_T_1 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 294:39]
  wire  _mem_WIRE_read_valid = 1'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire  _GEN_1960 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _GEN_1961 = _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:54]
  wire [5:0] _mem_WIRE_read_memWidth = 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [5:0] _GEN_1962 = 6'h8; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 290:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _GEN_1963 = 5'h0 == rd ? _next_reg_T_53 : _GEN_1743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1964 = 5'h1 == rd ? _next_reg_T_53 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1965 = 5'h2 == rd ? _next_reg_T_53 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1966 = 5'h3 == rd ? _next_reg_T_53 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1967 = 5'h4 == rd ? _next_reg_T_53 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1968 = 5'h5 == rd ? _next_reg_T_53 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1969 = 5'h6 == rd ? _next_reg_T_53 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1970 = 5'h7 == rd ? _next_reg_T_53 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1971 = 5'h8 == rd ? _next_reg_T_53 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1972 = 5'h9 == rd ? _next_reg_T_53 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1973 = 5'ha == rd ? _next_reg_T_53 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1974 = 5'hb == rd ? _next_reg_T_53 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1975 = 5'hc == rd ? _next_reg_T_53 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1976 = 5'hd == rd ? _next_reg_T_53 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1977 = 5'he == rd ? _next_reg_T_53 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1978 = 5'hf == rd ? _next_reg_T_53 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1979 = 5'h10 == rd ? _next_reg_T_53 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1980 = 5'h11 == rd ? _next_reg_T_53 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1981 = 5'h12 == rd ? _next_reg_T_53 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1982 = 5'h13 == rd ? _next_reg_T_53 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1983 = 5'h14 == rd ? _next_reg_T_53 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1984 = 5'h15 == rd ? _next_reg_T_53 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1985 = 5'h16 == rd ? _next_reg_T_53 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1986 = 5'h17 == rd ? _next_reg_T_53 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1987 = 5'h18 == rd ? _next_reg_T_53 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1988 = 5'h19 == rd ? _next_reg_T_53 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1989 = 5'h1a == rd ? _next_reg_T_53 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1990 = 5'h1b == rd ? _next_reg_T_53 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1991 = 5'h1c == rd ? _next_reg_T_53 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1992 = 5'h1d == rd ? _next_reg_T_53 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1993 = 5'h1e == rd ? _next_reg_T_53 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [31:0] _GEN_1994 = 5'h1f == rd ? _next_reg_T_53 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire  _GEN_1996 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [2:0] _GEN_2000 = _T_348 ? inst[14:12] : _GEN_1918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2002 = _T_348 ? inst[6:0] : _GEN_1921; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2004 = 32'h3 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _mem_WIRE_read_addr = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [31:0] _GEN_2005 = _T_348 ? _T_433 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [5:0] _GEN_2006 = _T_348 ? 6'h8 : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _GEN_2007 = _T_348 ? _GEN_1928 : _GEN_1743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2008 = _T_348 ? _GEN_1929 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2009 = _T_348 ? _GEN_1930 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2010 = _T_348 ? _GEN_1931 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2011 = _T_348 ? _GEN_1932 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2012 = _T_348 ? _GEN_1933 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2013 = _T_348 ? _GEN_1934 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2014 = _T_348 ? _GEN_1935 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2015 = _T_348 ? _GEN_1936 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2016 = _T_348 ? _GEN_1937 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2017 = _T_348 ? _GEN_1938 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2018 = _T_348 ? _GEN_1939 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2019 = _T_348 ? _GEN_1940 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2020 = _T_348 ? _GEN_1941 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2021 = _T_348 ? _GEN_1942 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2022 = _T_348 ? _GEN_1943 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2023 = _T_348 ? _GEN_1944 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2024 = _T_348 ? _GEN_1945 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2025 = _T_348 ? _GEN_1946 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2026 = _T_348 ? _GEN_1947 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2027 = _T_348 ? _GEN_1948 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2028 = _T_348 ? _GEN_1949 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2029 = _T_348 ? _GEN_1950 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2030 = _T_348 ? _GEN_1951 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2031 = _T_348 ? _GEN_1952 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2032 = _T_348 ? _GEN_1953 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2033 = _T_348 ? _GEN_1954 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2034 = _T_348 ? _GEN_1955 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2035 = _T_348 ? _GEN_1956 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2036 = _T_348 ? _GEN_1957 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2037 = _T_348 ? _GEN_1958 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [31:0] _GEN_2038 = _T_348 ? _GEN_1959 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire  _GEN_2040 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [2:0] _funct3_T_27 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_372 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_31 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_54 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:54]
  wire [31:0] _next_reg_T_55 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:54]
  wire [1:0] _next_reg_rOff_T_1 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_1 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_7 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_8 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_9 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_10 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_11 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_12 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_13 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_1 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_56 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_3341 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_57 = _GEN_3340 & 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [15:0] _next_reg_T_58 = _next_reg_T_57[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:66]
  wire  next_reg_signBit_1 = _next_reg_T_57[15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire  _next_reg_T_59 = next_reg_signBit_1; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [15:0] _next_reg_T_60 = next_reg_signBit_1 ? 16'hffff : 16'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [31:0] _next_reg_T_61 = {_next_reg_T_60,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _next_reg_rd_23 = {_next_reg_T_60,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [31:0] _GEN_2041 = 5'h0 == rd ? _next_reg_T_61 : _GEN_2007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2042 = 5'h1 == rd ? _next_reg_T_61 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2043 = 5'h2 == rd ? _next_reg_T_61 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2044 = 5'h3 == rd ? _next_reg_T_61 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2045 = 5'h4 == rd ? _next_reg_T_61 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2046 = 5'h5 == rd ? _next_reg_T_61 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2047 = 5'h6 == rd ? _next_reg_T_61 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2048 = 5'h7 == rd ? _next_reg_T_61 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2049 = 5'h8 == rd ? _next_reg_T_61 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2050 = 5'h9 == rd ? _next_reg_T_61 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2051 = 5'ha == rd ? _next_reg_T_61 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2052 = 5'hb == rd ? _next_reg_T_61 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2053 = 5'hc == rd ? _next_reg_T_61 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2054 = 5'hd == rd ? _next_reg_T_61 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2055 = 5'he == rd ? _next_reg_T_61 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2056 = 5'hf == rd ? _next_reg_T_61 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2057 = 5'h10 == rd ? _next_reg_T_61 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2058 = 5'h11 == rd ? _next_reg_T_61 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2059 = 5'h12 == rd ? _next_reg_T_61 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2060 = 5'h13 == rd ? _next_reg_T_61 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2061 = 5'h14 == rd ? _next_reg_T_61 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2062 = 5'h15 == rd ? _next_reg_T_61 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2063 = 5'h16 == rd ? _next_reg_T_61 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2064 = 5'h17 == rd ? _next_reg_T_61 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2065 = 5'h18 == rd ? _next_reg_T_61 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2066 = 5'h19 == rd ? _next_reg_T_61 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2067 = 5'h1a == rd ? _next_reg_T_61 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2068 = 5'h1b == rd ? _next_reg_T_61 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2069 = 5'h1c == rd ? _next_reg_T_61 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2070 = 5'h1d == rd ? _next_reg_T_61 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2071 = 5'h1e == rd ? _next_reg_T_61 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _GEN_2072 = 5'h1f == rd ? _next_reg_T_61 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [31:0] _now_reg_rs1_32 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 303:39]
  wire [31:0] _mem_read_addr_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 303:39]
  wire  _GEN_2073 = _T_435 | _T_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2074 = _T_435 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 303:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2075 = _T_435 ? 6'h10 : _GEN_2006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2076 = _T_435 ? _GEN_2041 : _GEN_2007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2077 = _T_435 ? _GEN_2042 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2078 = _T_435 ? _GEN_2043 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2079 = _T_435 ? _GEN_2044 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2080 = _T_435 ? _GEN_2045 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2081 = _T_435 ? _GEN_2046 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2082 = _T_435 ? _GEN_2047 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2083 = _T_435 ? _GEN_2048 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2084 = _T_435 ? _GEN_2049 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2085 = _T_435 ? _GEN_2050 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2086 = _T_435 ? _GEN_2051 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2087 = _T_435 ? _GEN_2052 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2088 = _T_435 ? _GEN_2053 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2089 = _T_435 ? _GEN_2054 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2090 = _T_435 ? _GEN_2055 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2091 = _T_435 ? _GEN_2056 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2092 = _T_435 ? _GEN_2057 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2093 = _T_435 ? _GEN_2058 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2094 = _T_435 ? _GEN_2059 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2095 = _T_435 ? _GEN_2060 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2096 = _T_435 ? _GEN_2061 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2097 = _T_435 ? _GEN_2062 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2098 = _T_435 ? _GEN_2063 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2099 = _T_435 ? _GEN_2064 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2100 = _T_435 ? _GEN_2065 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2101 = _T_435 ? _GEN_2066 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2102 = _T_435 ? _GEN_2067 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2103 = _T_435 ? _GEN_2068 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2104 = _T_435 ? _GEN_2069 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2105 = _T_435 ? _GEN_2070 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2106 = _T_435 ? _GEN_2071 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [31:0] _GEN_2107 = _T_435 ? _GEN_2072 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2109 = _T_435 ? _GEN_1926 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2113 = _T_368 ? inst[14:12] : _GEN_2000; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2115 = _T_368 ? inst[6:0] : _GEN_2002; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2117 = _T_368 ? _GEN_2073 : _T_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2118 = _T_368 ? _GEN_2074 : _GEN_2005; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [5:0] _GEN_2119 = _T_368 ? _GEN_2075 : _GEN_2006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2120 = _T_368 ? _GEN_2076 : _GEN_2007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2121 = _T_368 ? _GEN_2077 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2122 = _T_368 ? _GEN_2078 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2123 = _T_368 ? _GEN_2079 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2124 = _T_368 ? _GEN_2080 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2125 = _T_368 ? _GEN_2081 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2126 = _T_368 ? _GEN_2082 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2127 = _T_368 ? _GEN_2083 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2128 = _T_368 ? _GEN_2084 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2129 = _T_368 ? _GEN_2085 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2130 = _T_368 ? _GEN_2086 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2131 = _T_368 ? _GEN_2087 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2132 = _T_368 ? _GEN_2088 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2133 = _T_368 ? _GEN_2089 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2134 = _T_368 ? _GEN_2090 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2135 = _T_368 ? _GEN_2091 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2136 = _T_368 ? _GEN_2092 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2137 = _T_368 ? _GEN_2093 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2138 = _T_368 ? _GEN_2094 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2139 = _T_368 ? _GEN_2095 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2140 = _T_368 ? _GEN_2096 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2141 = _T_368 ? _GEN_2097 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2142 = _T_368 ? _GEN_2098 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2143 = _T_368 ? _GEN_2099 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2144 = _T_368 ? _GEN_2100 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2145 = _T_368 ? _GEN_2101 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2146 = _T_368 ? _GEN_2102 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2147 = _T_368 ? _GEN_2103 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2148 = _T_368 ? _GEN_2104 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2149 = _T_368 ? _GEN_2105 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2150 = _T_368 ? _GEN_2106 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [31:0] _GEN_2151 = _T_368 ? _GEN_2107 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2153 = _T_368 ? _GEN_2109 : _GEN_1926; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [2:0] _funct3_T_28 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_392 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_34 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_62 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:54]
  wire [31:0] _next_reg_T_63 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:54]
  wire [1:0] _next_reg_rOff_T_2 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_2 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_14 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_15 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_16 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_17 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_18 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_19 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_20 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_2 = 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_64 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_3342 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_65 = _GEN_3340 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [31:0] _next_reg_T_66 = _next_reg_T_65[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:66]
  wire  next_reg_signBit_2 = _next_reg_T_65[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_67 = _next_reg_T_65[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:66]
  wire [31:0] _next_reg_rd_24 = _next_reg_T_65[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:66]
  wire [31:0] _GEN_2154 = 5'h0 == rd ? _next_reg_T_65[31:0] : _GEN_2120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2155 = 5'h1 == rd ? _next_reg_T_65[31:0] : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2156 = 5'h2 == rd ? _next_reg_T_65[31:0] : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2157 = 5'h3 == rd ? _next_reg_T_65[31:0] : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2158 = 5'h4 == rd ? _next_reg_T_65[31:0] : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2159 = 5'h5 == rd ? _next_reg_T_65[31:0] : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2160 = 5'h6 == rd ? _next_reg_T_65[31:0] : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2161 = 5'h7 == rd ? _next_reg_T_65[31:0] : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2162 = 5'h8 == rd ? _next_reg_T_65[31:0] : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2163 = 5'h9 == rd ? _next_reg_T_65[31:0] : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2164 = 5'ha == rd ? _next_reg_T_65[31:0] : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2165 = 5'hb == rd ? _next_reg_T_65[31:0] : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2166 = 5'hc == rd ? _next_reg_T_65[31:0] : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2167 = 5'hd == rd ? _next_reg_T_65[31:0] : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2168 = 5'he == rd ? _next_reg_T_65[31:0] : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2169 = 5'hf == rd ? _next_reg_T_65[31:0] : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2170 = 5'h10 == rd ? _next_reg_T_65[31:0] : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2171 = 5'h11 == rd ? _next_reg_T_65[31:0] : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2172 = 5'h12 == rd ? _next_reg_T_65[31:0] : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2173 = 5'h13 == rd ? _next_reg_T_65[31:0] : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2174 = 5'h14 == rd ? _next_reg_T_65[31:0] : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2175 = 5'h15 == rd ? _next_reg_T_65[31:0] : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2176 = 5'h16 == rd ? _next_reg_T_65[31:0] : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2177 = 5'h17 == rd ? _next_reg_T_65[31:0] : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2178 = 5'h18 == rd ? _next_reg_T_65[31:0] : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2179 = 5'h19 == rd ? _next_reg_T_65[31:0] : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2180 = 5'h1a == rd ? _next_reg_T_65[31:0] : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2181 = 5'h1b == rd ? _next_reg_T_65[31:0] : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2182 = 5'h1c == rd ? _next_reg_T_65[31:0] : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2183 = 5'h1d == rd ? _next_reg_T_65[31:0] : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2184 = 5'h1e == rd ? _next_reg_T_65[31:0] : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _GEN_2185 = 5'h1f == rd ? _next_reg_T_65[31:0] : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [31:0] _now_reg_rs1_35 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T_4 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 312:39]
  wire [31:0] _mem_read_addr_T_5 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 312:39]
  wire  _GEN_2186 = _T_437 | _GEN_2117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2187 = _T_437 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 312:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2188 = _T_437 ? 6'h20 : _GEN_2119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2189 = _T_437 ? _GEN_2154 : _GEN_2120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2190 = _T_437 ? _GEN_2155 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2191 = _T_437 ? _GEN_2156 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2192 = _T_437 ? _GEN_2157 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2193 = _T_437 ? _GEN_2158 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2194 = _T_437 ? _GEN_2159 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2195 = _T_437 ? _GEN_2160 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2196 = _T_437 ? _GEN_2161 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2197 = _T_437 ? _GEN_2162 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2198 = _T_437 ? _GEN_2163 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2199 = _T_437 ? _GEN_2164 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2200 = _T_437 ? _GEN_2165 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2201 = _T_437 ? _GEN_2166 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2202 = _T_437 ? _GEN_2167 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2203 = _T_437 ? _GEN_2168 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2204 = _T_437 ? _GEN_2169 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2205 = _T_437 ? _GEN_2170 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2206 = _T_437 ? _GEN_2171 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2207 = _T_437 ? _GEN_2172 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2208 = _T_437 ? _GEN_2173 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2209 = _T_437 ? _GEN_2174 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2210 = _T_437 ? _GEN_2175 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2211 = _T_437 ? _GEN_2176 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2212 = _T_437 ? _GEN_2177 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2213 = _T_437 ? _GEN_2178 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2214 = _T_437 ? _GEN_2179 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2215 = _T_437 ? _GEN_2180 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2216 = _T_437 ? _GEN_2181 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2217 = _T_437 ? _GEN_2182 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2218 = _T_437 ? _GEN_2183 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2219 = _T_437 ? _GEN_2184 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [31:0] _GEN_2220 = _T_437 ? _GEN_2185 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2222 = _T_437 ? _GEN_2153 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2226 = _T_388 ? inst[14:12] : _GEN_2113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2228 = _T_388 ? inst[6:0] : _GEN_2115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2230 = _T_388 ? _GEN_2186 : _GEN_2117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2231 = _T_388 ? _GEN_2187 : _GEN_2118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [5:0] _GEN_2232 = _T_388 ? _GEN_2188 : _GEN_2119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2233 = _T_388 ? _GEN_2189 : _GEN_2120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2234 = _T_388 ? _GEN_2190 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2235 = _T_388 ? _GEN_2191 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2236 = _T_388 ? _GEN_2192 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2237 = _T_388 ? _GEN_2193 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2238 = _T_388 ? _GEN_2194 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2239 = _T_388 ? _GEN_2195 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2240 = _T_388 ? _GEN_2196 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2241 = _T_388 ? _GEN_2197 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2242 = _T_388 ? _GEN_2198 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2243 = _T_388 ? _GEN_2199 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2244 = _T_388 ? _GEN_2200 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2245 = _T_388 ? _GEN_2201 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2246 = _T_388 ? _GEN_2202 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2247 = _T_388 ? _GEN_2203 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2248 = _T_388 ? _GEN_2204 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2249 = _T_388 ? _GEN_2205 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2250 = _T_388 ? _GEN_2206 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2251 = _T_388 ? _GEN_2207 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2252 = _T_388 ? _GEN_2208 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2253 = _T_388 ? _GEN_2209 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2254 = _T_388 ? _GEN_2210 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2255 = _T_388 ? _GEN_2211 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2256 = _T_388 ? _GEN_2212 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2257 = _T_388 ? _GEN_2213 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2258 = _T_388 ? _GEN_2214 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2259 = _T_388 ? _GEN_2215 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2260 = _T_388 ? _GEN_2216 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2261 = _T_388 ? _GEN_2217 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2262 = _T_388 ? _GEN_2218 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2263 = _T_388 ? _GEN_2219 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _GEN_2264 = _T_388 ? _GEN_2220 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2266 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [2:0] _funct3_T_29 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_412 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _GEN_2268 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [31:0] _now_reg_rs1_36 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_68 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:118]
  wire [31:0] _next_reg_T_69 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:118]
  wire [1:0] _next_reg_rOff_T_3 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_3 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_21 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_22 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_23 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_24 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_25 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_26 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_27 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_3 = 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_70 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_3343 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_71 = _GEN_3340 & 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [7:0] _next_reg_T_72 = _next_reg_T_49[7:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:129]
  wire [31:0] _next_reg_T_73 = {24'h0,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_reg_rd_25 = {24'h0,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_2269 = 5'h0 == rd ? _next_reg_T_73 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2270 = 5'h1 == rd ? _next_reg_T_73 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2271 = 5'h2 == rd ? _next_reg_T_73 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2272 = 5'h3 == rd ? _next_reg_T_73 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2273 = 5'h4 == rd ? _next_reg_T_73 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2274 = 5'h5 == rd ? _next_reg_T_73 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2275 = 5'h6 == rd ? _next_reg_T_73 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2276 = 5'h7 == rd ? _next_reg_T_73 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2277 = 5'h8 == rd ? _next_reg_T_73 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2278 = 5'h9 == rd ? _next_reg_T_73 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2279 = 5'ha == rd ? _next_reg_T_73 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2280 = 5'hb == rd ? _next_reg_T_73 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2281 = 5'hc == rd ? _next_reg_T_73 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2282 = 5'hd == rd ? _next_reg_T_73 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2283 = 5'he == rd ? _next_reg_T_73 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2284 = 5'hf == rd ? _next_reg_T_73 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2285 = 5'h10 == rd ? _next_reg_T_73 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2286 = 5'h11 == rd ? _next_reg_T_73 : _GEN_2250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2287 = 5'h12 == rd ? _next_reg_T_73 : _GEN_2251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2288 = 5'h13 == rd ? _next_reg_T_73 : _GEN_2252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2289 = 5'h14 == rd ? _next_reg_T_73 : _GEN_2253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2290 = 5'h15 == rd ? _next_reg_T_73 : _GEN_2254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2291 = 5'h16 == rd ? _next_reg_T_73 : _GEN_2255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2292 = 5'h17 == rd ? _next_reg_T_73 : _GEN_2256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2293 = 5'h18 == rd ? _next_reg_T_73 : _GEN_2257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2294 = 5'h19 == rd ? _next_reg_T_73 : _GEN_2258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2295 = 5'h1a == rd ? _next_reg_T_73 : _GEN_2259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2296 = 5'h1b == rd ? _next_reg_T_73 : _GEN_2260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2297 = 5'h1c == rd ? _next_reg_T_73 : _GEN_2261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2298 = 5'h1d == rd ? _next_reg_T_73 : _GEN_2262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2299 = 5'h1e == rd ? _next_reg_T_73 : _GEN_2263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [31:0] _GEN_2300 = 5'h1f == rd ? _next_reg_T_73 : _GEN_2264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [2:0] _GEN_2304 = _T_408 ? inst[14:12] : _GEN_2226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2306 = _T_408 ? inst[6:0] : _GEN_2228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2309 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2310 = _T_408 | _GEN_2230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2311 = _T_408 ? _T_433 : _GEN_2231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2312 = _T_408 ? 6'h8 : _GEN_2232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2313 = _T_408 ? _GEN_2269 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2314 = _T_408 ? _GEN_2270 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2315 = _T_408 ? _GEN_2271 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2316 = _T_408 ? _GEN_2272 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2317 = _T_408 ? _GEN_2273 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2318 = _T_408 ? _GEN_2274 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2319 = _T_408 ? _GEN_2275 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2320 = _T_408 ? _GEN_2276 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2321 = _T_408 ? _GEN_2277 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2322 = _T_408 ? _GEN_2278 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2323 = _T_408 ? _GEN_2279 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2324 = _T_408 ? _GEN_2280 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2325 = _T_408 ? _GEN_2281 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2326 = _T_408 ? _GEN_2282 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2327 = _T_408 ? _GEN_2283 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2328 = _T_408 ? _GEN_2284 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2329 = _T_408 ? _GEN_2285 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2330 = _T_408 ? _GEN_2286 : _GEN_2250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2331 = _T_408 ? _GEN_2287 : _GEN_2251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2332 = _T_408 ? _GEN_2288 : _GEN_2252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2333 = _T_408 ? _GEN_2289 : _GEN_2253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2334 = _T_408 ? _GEN_2290 : _GEN_2254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2335 = _T_408 ? _GEN_2291 : _GEN_2255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2336 = _T_408 ? _GEN_2292 : _GEN_2256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2337 = _T_408 ? _GEN_2293 : _GEN_2257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2338 = _T_408 ? _GEN_2294 : _GEN_2258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2339 = _T_408 ? _GEN_2295 : _GEN_2259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2340 = _T_408 ? _GEN_2296 : _GEN_2260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2341 = _T_408 ? _GEN_2297 : _GEN_2261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2342 = _T_408 ? _GEN_2298 : _GEN_2262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2343 = _T_408 ? _GEN_2299 : _GEN_2263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [31:0] _GEN_2344 = _T_408 ? _GEN_2300 : _GEN_2264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [2:0] _funct3_T_30 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_431 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_38 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _next_reg_T_74 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:54]
  wire [31:0] _next_reg_T_75 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:54]
  wire [1:0] _next_reg_rOff_T_4 = _T_433[1:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:28]
  wire [4:0] next_reg_rOff_4 = {_T_433[1:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire  _next_reg_rMask_T_28 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_29 = 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_30 = 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_31 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_32 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] _next_reg_rMask_T_33 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire  _next_reg_rMask_T_34 = 1'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [63:0] next_reg_rMask_4 = 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 38:32]
  wire [31:0] _next_reg_T_76 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _GEN_3344 = {{32'd0}, _next_reg_T_48}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [63:0] _next_reg_T_77 = _GEN_3340 & 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire [15:0] _next_reg_T_78 = _next_reg_T_57[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:66]
  wire [31:0] _next_reg_T_79 = {16'h0,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_reg_rd_26 = {16'h0,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_2345 = 5'h0 == rd ? _next_reg_T_79 : _GEN_2313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2346 = 5'h1 == rd ? _next_reg_T_79 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2347 = 5'h2 == rd ? _next_reg_T_79 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2348 = 5'h3 == rd ? _next_reg_T_79 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2349 = 5'h4 == rd ? _next_reg_T_79 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2350 = 5'h5 == rd ? _next_reg_T_79 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2351 = 5'h6 == rd ? _next_reg_T_79 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2352 = 5'h7 == rd ? _next_reg_T_79 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2353 = 5'h8 == rd ? _next_reg_T_79 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2354 = 5'h9 == rd ? _next_reg_T_79 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2355 = 5'ha == rd ? _next_reg_T_79 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2356 = 5'hb == rd ? _next_reg_T_79 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2357 = 5'hc == rd ? _next_reg_T_79 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2358 = 5'hd == rd ? _next_reg_T_79 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2359 = 5'he == rd ? _next_reg_T_79 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2360 = 5'hf == rd ? _next_reg_T_79 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2361 = 5'h10 == rd ? _next_reg_T_79 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2362 = 5'h11 == rd ? _next_reg_T_79 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2363 = 5'h12 == rd ? _next_reg_T_79 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2364 = 5'h13 == rd ? _next_reg_T_79 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2365 = 5'h14 == rd ? _next_reg_T_79 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2366 = 5'h15 == rd ? _next_reg_T_79 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2367 = 5'h16 == rd ? _next_reg_T_79 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2368 = 5'h17 == rd ? _next_reg_T_79 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2369 = 5'h18 == rd ? _next_reg_T_79 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2370 = 5'h19 == rd ? _next_reg_T_79 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2371 = 5'h1a == rd ? _next_reg_T_79 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2372 = 5'h1b == rd ? _next_reg_T_79 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2373 = 5'h1c == rd ? _next_reg_T_79 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2374 = 5'h1d == rd ? _next_reg_T_79 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2375 = 5'h1e == rd ? _next_reg_T_79 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _GEN_2376 = 5'h1f == rd ? _next_reg_T_79 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [31:0] _now_reg_rs1_39 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_read_addr_T_6 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 322:39]
  wire [31:0] _mem_read_addr_T_7 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 322:39]
  wire  _GEN_2377 = _T_435 | _GEN_2310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [31:0] _GEN_2378 = _T_435 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 322:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [5:0] _GEN_2379 = _T_435 ? 6'h10 : _GEN_2312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [31:0] _GEN_2380 = _T_435 ? _GEN_2345 : _GEN_2313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2381 = _T_435 ? _GEN_2346 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2382 = _T_435 ? _GEN_2347 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2383 = _T_435 ? _GEN_2348 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2384 = _T_435 ? _GEN_2349 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2385 = _T_435 ? _GEN_2350 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2386 = _T_435 ? _GEN_2351 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2387 = _T_435 ? _GEN_2352 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2388 = _T_435 ? _GEN_2353 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2389 = _T_435 ? _GEN_2354 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2390 = _T_435 ? _GEN_2355 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2391 = _T_435 ? _GEN_2356 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2392 = _T_435 ? _GEN_2357 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2393 = _T_435 ? _GEN_2358 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2394 = _T_435 ? _GEN_2359 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2395 = _T_435 ? _GEN_2360 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2396 = _T_435 ? _GEN_2361 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2397 = _T_435 ? _GEN_2362 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2398 = _T_435 ? _GEN_2363 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2399 = _T_435 ? _GEN_2364 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2400 = _T_435 ? _GEN_2365 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2401 = _T_435 ? _GEN_2366 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2402 = _T_435 ? _GEN_2367 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2403 = _T_435 ? _GEN_2368 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2404 = _T_435 ? _GEN_2369 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2405 = _T_435 ? _GEN_2370 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2406 = _T_435 ? _GEN_2371 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2407 = _T_435 ? _GEN_2372 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2408 = _T_435 ? _GEN_2373 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2409 = _T_435 ? _GEN_2374 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2410 = _T_435 ? _GEN_2375 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [31:0] _GEN_2411 = _T_435 ? _GEN_2376 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_2413 = _T_435 ? _GEN_2266 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2417 = _T_427 ? inst[14:12] : _GEN_2304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2419 = _T_427 ? inst[6:0] : _GEN_2306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2421 = _T_427 ? _GEN_2377 : _GEN_2310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2422 = _T_427 ? _GEN_2074 : _GEN_2311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [5:0] _GEN_2423 = _T_427 ? _GEN_2379 : _GEN_2312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2424 = _T_427 ? _GEN_2380 : _GEN_2313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2425 = _T_427 ? _GEN_2381 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2426 = _T_427 ? _GEN_2382 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2427 = _T_427 ? _GEN_2383 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2428 = _T_427 ? _GEN_2384 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2429 = _T_427 ? _GEN_2385 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2430 = _T_427 ? _GEN_2386 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2431 = _T_427 ? _GEN_2387 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2432 = _T_427 ? _GEN_2388 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2433 = _T_427 ? _GEN_2389 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2434 = _T_427 ? _GEN_2390 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2435 = _T_427 ? _GEN_2391 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2436 = _T_427 ? _GEN_2392 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2437 = _T_427 ? _GEN_2393 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2438 = _T_427 ? _GEN_2394 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2439 = _T_427 ? _GEN_2395 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2440 = _T_427 ? _GEN_2396 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2441 = _T_427 ? _GEN_2397 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2442 = _T_427 ? _GEN_2398 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2443 = _T_427 ? _GEN_2399 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2444 = _T_427 ? _GEN_2400 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2445 = _T_427 ? _GEN_2401 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2446 = _T_427 ? _GEN_2402 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2447 = _T_427 ? _GEN_2403 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2448 = _T_427 ? _GEN_2404 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2449 = _T_427 ? _GEN_2405 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2450 = _T_427 ? _GEN_2406 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2451 = _T_427 ? _GEN_2407 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2452 = _T_427 ? _GEN_2408 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2453 = _T_427 ? _GEN_2409 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2454 = _T_427 ? _GEN_2410 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _GEN_2455 = _T_427 ? _GEN_2411 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_2457 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [2:0] _funct3_T_31 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_452 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _GEN_2459 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [31:0] _now_reg_rs1_40 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_466 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:95]
  wire [31:0] _T_467 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:95]
  wire [31:0] _now_reg_rs2_15 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [7:0] _T_468 = _GEN_840[7:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:119]
  wire [2:0] _GEN_2464 = _T_447 ? inst[14:12] : _GEN_2417; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2466 = _T_447 ? inst[6:0] : _GEN_2419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2469 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _mem_WIRE_write_valid = 1'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire  _GEN_2470 = 32'h23 == _T_426; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _mem_WIRE_write_addr = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [31:0] _GEN_2471 = _T_447 ? _T_433 : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [5:0] _mem_WIRE_write_memWidth = 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [5:0] _GEN_2472 = _T_447 ? 6'h8 : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [31:0] _mem_WIRE_write_data = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire [31:0] _GEN_2473 = _T_447 ? {{24'd0}, _GEN_840[7:0]} : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [2:0] _funct3_T_32 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_475 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_42 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_490 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 331:31]
  wire [31:0] _T_491 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 331:31]
  wire [31:0] _now_reg_rs2_16 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [15:0] _T_492 = _GEN_840[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 331:56]
  wire [31:0] _now_reg_rs1_43 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_write_addr_T = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 333:40]
  wire [31:0] _mem_write_addr_T_1 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 333:40]
  wire  _GEN_2474 = _T_435 | _T_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [31:0] _GEN_2475 = _T_435 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 333:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [5:0] _GEN_2476 = _T_435 ? 6'h10 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [31:0] _GEN_2477 = _T_435 ? {{16'd0}, _GEN_840[15:0]} : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_2479 = _T_435 ? _GEN_2457 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2484 = _T_470 ? inst[14:12] : _GEN_2464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2486 = _T_470 ? inst[6:0] : _GEN_2466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2488 = _T_470 ? _GEN_2474 : _T_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [31:0] _GEN_2489 = _T_470 ? _GEN_2074 : _GEN_2471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [5:0] _GEN_2490 = _T_470 ? _GEN_2476 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [31:0] _GEN_2491 = _T_470 ? _GEN_2477 : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2493 = _T_470 ? _GEN_2479 : _GEN_2457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [2:0] _funct3_T_33 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_499 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_45 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _T_514 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 340:31]
  wire [31:0] _T_515 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 340:31]
  wire [31:0] _now_reg_rs2_17 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _T_516 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _now_reg_rs1_46 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [32:0] _mem_write_addr_T_2 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 342:40]
  wire [31:0] _mem_write_addr_T_3 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 342:40]
  wire  _GEN_2494 = _T_437 | _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [31:0] _GEN_2495 = _T_437 ? _T_433 : _T_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 342:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [5:0] _GEN_2496 = _T_437 ? 6'h20 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [31:0] _GEN_2497 = _T_437 ? _GEN_840 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_2499 = _T_437 ? _GEN_2493 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2504 = _T_494 ? inst[14:12] : _GEN_2484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2506 = _T_494 ? inst[6:0] : _GEN_2486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2508 = _T_494 ? _GEN_2494 : _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [31:0] _GEN_2509 = _T_494 ? _GEN_2187 : _GEN_2489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [5:0] _GEN_2510 = _T_494 ? _GEN_2496 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [31:0] _GEN_2511 = _T_494 ? _GEN_2497 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_2513 = _T_494 ? _GEN_2499 : _GEN_2493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [2:0] _funct3_T_34 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_522 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_2517 = _T_518 ? inst[14:12] : _GEN_2504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2519 = _T_518 ? inst[6:0] : _GEN_2506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2522 = _T_518 | _GEN_2513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _funct3_T_35 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_528 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  _GEN_2524 = 2'h0 == io_now_internal_privilegeMode | _GEN_2522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2526 = 2'h1 == io_now_internal_privilegeMode | (2'h0 == io_now_internal_privilegeMode | _GEN_2522); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2529 = 2'h3 == io_now_internal_privilegeMode | (2'h1 == io_now_internal_privilegeMode | (2'h0 ==
    io_now_internal_privilegeMode | _GEN_2522)); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [2:0] _GEN_2535 = _T_524 ? inst[14:12] : _GEN_2517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2537 = _T_524 ? inst[6:0] : _GEN_2519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire  _GEN_2540 = _T_524 ? _GEN_2529 : _GEN_2522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23]
  wire [2:0] _funct3_T_36 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_537 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_2546 = _T_533 ? inst[14:12] : _GEN_2535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2548 = _T_533 ? inst[6:0] : _GEN_2537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [6:0] _funct7_T_10 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_37 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_544 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_47 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_18 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _next_reg_T_80 = _GEN_31 * _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:65]
  wire [31:0] _next_reg_T_81 = _next_reg_T_80[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:80]
  wire [31:0] _next_reg_rd_27 = _next_reg_T_80[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:80]
  wire [31:0] _GEN_2550 = 5'h0 == rd ? _next_reg_T_80[31:0] : _GEN_2424; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2551 = 5'h1 == rd ? _next_reg_T_80[31:0] : _GEN_2425; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2552 = 5'h2 == rd ? _next_reg_T_80[31:0] : _GEN_2426; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2553 = 5'h3 == rd ? _next_reg_T_80[31:0] : _GEN_2427; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2554 = 5'h4 == rd ? _next_reg_T_80[31:0] : _GEN_2428; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2555 = 5'h5 == rd ? _next_reg_T_80[31:0] : _GEN_2429; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2556 = 5'h6 == rd ? _next_reg_T_80[31:0] : _GEN_2430; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2557 = 5'h7 == rd ? _next_reg_T_80[31:0] : _GEN_2431; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2558 = 5'h8 == rd ? _next_reg_T_80[31:0] : _GEN_2432; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2559 = 5'h9 == rd ? _next_reg_T_80[31:0] : _GEN_2433; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2560 = 5'ha == rd ? _next_reg_T_80[31:0] : _GEN_2434; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2561 = 5'hb == rd ? _next_reg_T_80[31:0] : _GEN_2435; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2562 = 5'hc == rd ? _next_reg_T_80[31:0] : _GEN_2436; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2563 = 5'hd == rd ? _next_reg_T_80[31:0] : _GEN_2437; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2564 = 5'he == rd ? _next_reg_T_80[31:0] : _GEN_2438; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2565 = 5'hf == rd ? _next_reg_T_80[31:0] : _GEN_2439; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2566 = 5'h10 == rd ? _next_reg_T_80[31:0] : _GEN_2440; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2567 = 5'h11 == rd ? _next_reg_T_80[31:0] : _GEN_2441; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2568 = 5'h12 == rd ? _next_reg_T_80[31:0] : _GEN_2442; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2569 = 5'h13 == rd ? _next_reg_T_80[31:0] : _GEN_2443; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2570 = 5'h14 == rd ? _next_reg_T_80[31:0] : _GEN_2444; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2571 = 5'h15 == rd ? _next_reg_T_80[31:0] : _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2572 = 5'h16 == rd ? _next_reg_T_80[31:0] : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2573 = 5'h17 == rd ? _next_reg_T_80[31:0] : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2574 = 5'h18 == rd ? _next_reg_T_80[31:0] : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2575 = 5'h19 == rd ? _next_reg_T_80[31:0] : _GEN_2449; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2576 = 5'h1a == rd ? _next_reg_T_80[31:0] : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2577 = 5'h1b == rd ? _next_reg_T_80[31:0] : _GEN_2451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2578 = 5'h1c == rd ? _next_reg_T_80[31:0] : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2579 = 5'h1d == rd ? _next_reg_T_80[31:0] : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2580 = 5'h1e == rd ? _next_reg_T_80[31:0] : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [31:0] _GEN_2581 = 5'h1f == rd ? _next_reg_T_80[31:0] : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [6:0] _GEN_2583 = _T_539 ? inst[31:25] : _GEN_1513; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2586 = _T_539 ? inst[14:12] : _GEN_2546; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2588 = _T_539 ? inst[6:0] : _GEN_2548; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2589 = _T_539 ? _GEN_2550 : _GEN_2424; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2590 = _T_539 ? _GEN_2551 : _GEN_2425; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2591 = _T_539 ? _GEN_2552 : _GEN_2426; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2592 = _T_539 ? _GEN_2553 : _GEN_2427; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2593 = _T_539 ? _GEN_2554 : _GEN_2428; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2594 = _T_539 ? _GEN_2555 : _GEN_2429; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2595 = _T_539 ? _GEN_2556 : _GEN_2430; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2596 = _T_539 ? _GEN_2557 : _GEN_2431; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2597 = _T_539 ? _GEN_2558 : _GEN_2432; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2598 = _T_539 ? _GEN_2559 : _GEN_2433; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2599 = _T_539 ? _GEN_2560 : _GEN_2434; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2600 = _T_539 ? _GEN_2561 : _GEN_2435; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2601 = _T_539 ? _GEN_2562 : _GEN_2436; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2602 = _T_539 ? _GEN_2563 : _GEN_2437; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2603 = _T_539 ? _GEN_2564 : _GEN_2438; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2604 = _T_539 ? _GEN_2565 : _GEN_2439; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2605 = _T_539 ? _GEN_2566 : _GEN_2440; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2606 = _T_539 ? _GEN_2567 : _GEN_2441; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2607 = _T_539 ? _GEN_2568 : _GEN_2442; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2608 = _T_539 ? _GEN_2569 : _GEN_2443; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2609 = _T_539 ? _GEN_2570 : _GEN_2444; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2610 = _T_539 ? _GEN_2571 : _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2611 = _T_539 ? _GEN_2572 : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2612 = _T_539 ? _GEN_2573 : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2613 = _T_539 ? _GEN_2574 : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2614 = _T_539 ? _GEN_2575 : _GEN_2449; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2615 = _T_539 ? _GEN_2576 : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2616 = _T_539 ? _GEN_2577 : _GEN_2451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2617 = _T_539 ? _GEN_2578 : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2618 = _T_539 ? _GEN_2579 : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2619 = _T_539 ? _GEN_2580 : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [31:0] _GEN_2620 = _T_539 ? _GEN_2581 : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [6:0] _funct7_T_11 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_38 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_551 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_48 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_82 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:65]
  wire [31:0] _now_reg_rs2_19 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_83 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:87]
  wire [63:0] _next_reg_T_84 = $signed(_T_300) * $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:72]
  wire [63:0] _next_reg_T_85 = $signed(_T_300) * $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:95]
  wire [31:0] _next_reg_T_86 = _next_reg_T_85[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:101]
  wire [31:0] _next_reg_rd_28 = _next_reg_T_85[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:101]
  wire [31:0] _GEN_2621 = 5'h0 == rd ? _next_reg_T_85[63:32] : _GEN_2589; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2622 = 5'h1 == rd ? _next_reg_T_85[63:32] : _GEN_2590; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2623 = 5'h2 == rd ? _next_reg_T_85[63:32] : _GEN_2591; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2624 = 5'h3 == rd ? _next_reg_T_85[63:32] : _GEN_2592; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2625 = 5'h4 == rd ? _next_reg_T_85[63:32] : _GEN_2593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2626 = 5'h5 == rd ? _next_reg_T_85[63:32] : _GEN_2594; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2627 = 5'h6 == rd ? _next_reg_T_85[63:32] : _GEN_2595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2628 = 5'h7 == rd ? _next_reg_T_85[63:32] : _GEN_2596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2629 = 5'h8 == rd ? _next_reg_T_85[63:32] : _GEN_2597; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2630 = 5'h9 == rd ? _next_reg_T_85[63:32] : _GEN_2598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2631 = 5'ha == rd ? _next_reg_T_85[63:32] : _GEN_2599; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2632 = 5'hb == rd ? _next_reg_T_85[63:32] : _GEN_2600; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2633 = 5'hc == rd ? _next_reg_T_85[63:32] : _GEN_2601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2634 = 5'hd == rd ? _next_reg_T_85[63:32] : _GEN_2602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2635 = 5'he == rd ? _next_reg_T_85[63:32] : _GEN_2603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2636 = 5'hf == rd ? _next_reg_T_85[63:32] : _GEN_2604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2637 = 5'h10 == rd ? _next_reg_T_85[63:32] : _GEN_2605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2638 = 5'h11 == rd ? _next_reg_T_85[63:32] : _GEN_2606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2639 = 5'h12 == rd ? _next_reg_T_85[63:32] : _GEN_2607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2640 = 5'h13 == rd ? _next_reg_T_85[63:32] : _GEN_2608; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2641 = 5'h14 == rd ? _next_reg_T_85[63:32] : _GEN_2609; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2642 = 5'h15 == rd ? _next_reg_T_85[63:32] : _GEN_2610; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2643 = 5'h16 == rd ? _next_reg_T_85[63:32] : _GEN_2611; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2644 = 5'h17 == rd ? _next_reg_T_85[63:32] : _GEN_2612; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2645 = 5'h18 == rd ? _next_reg_T_85[63:32] : _GEN_2613; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2646 = 5'h19 == rd ? _next_reg_T_85[63:32] : _GEN_2614; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2647 = 5'h1a == rd ? _next_reg_T_85[63:32] : _GEN_2615; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2648 = 5'h1b == rd ? _next_reg_T_85[63:32] : _GEN_2616; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2649 = 5'h1c == rd ? _next_reg_T_85[63:32] : _GEN_2617; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2650 = 5'h1d == rd ? _next_reg_T_85[63:32] : _GEN_2618; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2651 = 5'h1e == rd ? _next_reg_T_85[63:32] : _GEN_2619; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [31:0] _GEN_2652 = 5'h1f == rd ? _next_reg_T_85[63:32] : _GEN_2620; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [6:0] _GEN_2654 = _T_546 ? inst[31:25] : _GEN_2583; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2657 = _T_546 ? inst[14:12] : _GEN_2586; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2659 = _T_546 ? inst[6:0] : _GEN_2588; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2660 = _T_546 ? _GEN_2621 : _GEN_2589; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2661 = _T_546 ? _GEN_2622 : _GEN_2590; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2662 = _T_546 ? _GEN_2623 : _GEN_2591; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2663 = _T_546 ? _GEN_2624 : _GEN_2592; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2664 = _T_546 ? _GEN_2625 : _GEN_2593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2665 = _T_546 ? _GEN_2626 : _GEN_2594; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2666 = _T_546 ? _GEN_2627 : _GEN_2595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2667 = _T_546 ? _GEN_2628 : _GEN_2596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2668 = _T_546 ? _GEN_2629 : _GEN_2597; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2669 = _T_546 ? _GEN_2630 : _GEN_2598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2670 = _T_546 ? _GEN_2631 : _GEN_2599; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2671 = _T_546 ? _GEN_2632 : _GEN_2600; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2672 = _T_546 ? _GEN_2633 : _GEN_2601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2673 = _T_546 ? _GEN_2634 : _GEN_2602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2674 = _T_546 ? _GEN_2635 : _GEN_2603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2675 = _T_546 ? _GEN_2636 : _GEN_2604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2676 = _T_546 ? _GEN_2637 : _GEN_2605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2677 = _T_546 ? _GEN_2638 : _GEN_2606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2678 = _T_546 ? _GEN_2639 : _GEN_2607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2679 = _T_546 ? _GEN_2640 : _GEN_2608; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2680 = _T_546 ? _GEN_2641 : _GEN_2609; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2681 = _T_546 ? _GEN_2642 : _GEN_2610; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2682 = _T_546 ? _GEN_2643 : _GEN_2611; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2683 = _T_546 ? _GEN_2644 : _GEN_2612; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2684 = _T_546 ? _GEN_2645 : _GEN_2613; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2685 = _T_546 ? _GEN_2646 : _GEN_2614; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2686 = _T_546 ? _GEN_2647 : _GEN_2615; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2687 = _T_546 ? _GEN_2648 : _GEN_2616; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2688 = _T_546 ? _GEN_2649 : _GEN_2617; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2689 = _T_546 ? _GEN_2650 : _GEN_2618; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2690 = _T_546 ? _GEN_2651 : _GEN_2619; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [31:0] _GEN_2691 = _T_546 ? _GEN_2652 : _GEN_2620; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [6:0] _funct7_T_12 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_39 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_558 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_49 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_87 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:65]
  wire [31:0] _now_reg_rs2_20 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [32:0] _next_reg_T_88 = {1'b0,$signed(_GEN_840)}; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [64:0] _next_reg_T_89 = $signed(_T_300) * $signed(_next_reg_T_88); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [63:0] _next_reg_T_90 = _next_reg_T_89[63:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [63:0] _next_reg_T_91 = _next_reg_T_89[63:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [63:0] _next_reg_T_92 = _next_reg_T_89[63:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:88]
  wire [31:0] _next_reg_T_93 = _next_reg_T_92[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:94]
  wire [31:0] _next_reg_rd_29 = _next_reg_T_92[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:94]
  wire [31:0] _GEN_2692 = 5'h0 == rd ? _next_reg_T_92[63:32] : _GEN_2660; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2693 = 5'h1 == rd ? _next_reg_T_92[63:32] : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2694 = 5'h2 == rd ? _next_reg_T_92[63:32] : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2695 = 5'h3 == rd ? _next_reg_T_92[63:32] : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2696 = 5'h4 == rd ? _next_reg_T_92[63:32] : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2697 = 5'h5 == rd ? _next_reg_T_92[63:32] : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2698 = 5'h6 == rd ? _next_reg_T_92[63:32] : _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2699 = 5'h7 == rd ? _next_reg_T_92[63:32] : _GEN_2667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2700 = 5'h8 == rd ? _next_reg_T_92[63:32] : _GEN_2668; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2701 = 5'h9 == rd ? _next_reg_T_92[63:32] : _GEN_2669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2702 = 5'ha == rd ? _next_reg_T_92[63:32] : _GEN_2670; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2703 = 5'hb == rd ? _next_reg_T_92[63:32] : _GEN_2671; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2704 = 5'hc == rd ? _next_reg_T_92[63:32] : _GEN_2672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2705 = 5'hd == rd ? _next_reg_T_92[63:32] : _GEN_2673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2706 = 5'he == rd ? _next_reg_T_92[63:32] : _GEN_2674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2707 = 5'hf == rd ? _next_reg_T_92[63:32] : _GEN_2675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2708 = 5'h10 == rd ? _next_reg_T_92[63:32] : _GEN_2676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2709 = 5'h11 == rd ? _next_reg_T_92[63:32] : _GEN_2677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2710 = 5'h12 == rd ? _next_reg_T_92[63:32] : _GEN_2678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2711 = 5'h13 == rd ? _next_reg_T_92[63:32] : _GEN_2679; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2712 = 5'h14 == rd ? _next_reg_T_92[63:32] : _GEN_2680; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2713 = 5'h15 == rd ? _next_reg_T_92[63:32] : _GEN_2681; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2714 = 5'h16 == rd ? _next_reg_T_92[63:32] : _GEN_2682; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2715 = 5'h17 == rd ? _next_reg_T_92[63:32] : _GEN_2683; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2716 = 5'h18 == rd ? _next_reg_T_92[63:32] : _GEN_2684; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2717 = 5'h19 == rd ? _next_reg_T_92[63:32] : _GEN_2685; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2718 = 5'h1a == rd ? _next_reg_T_92[63:32] : _GEN_2686; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2719 = 5'h1b == rd ? _next_reg_T_92[63:32] : _GEN_2687; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2720 = 5'h1c == rd ? _next_reg_T_92[63:32] : _GEN_2688; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2721 = 5'h1d == rd ? _next_reg_T_92[63:32] : _GEN_2689; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2722 = 5'h1e == rd ? _next_reg_T_92[63:32] : _GEN_2690; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [31:0] _GEN_2723 = 5'h1f == rd ? _next_reg_T_92[63:32] : _GEN_2691; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [6:0] _GEN_2725 = _T_553 ? inst[31:25] : _GEN_2654; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2728 = _T_553 ? inst[14:12] : _GEN_2657; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2730 = _T_553 ? inst[6:0] : _GEN_2659; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2731 = _T_553 ? _GEN_2692 : _GEN_2660; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2732 = _T_553 ? _GEN_2693 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2733 = _T_553 ? _GEN_2694 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2734 = _T_553 ? _GEN_2695 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2735 = _T_553 ? _GEN_2696 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2736 = _T_553 ? _GEN_2697 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2737 = _T_553 ? _GEN_2698 : _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2738 = _T_553 ? _GEN_2699 : _GEN_2667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2739 = _T_553 ? _GEN_2700 : _GEN_2668; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2740 = _T_553 ? _GEN_2701 : _GEN_2669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2741 = _T_553 ? _GEN_2702 : _GEN_2670; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2742 = _T_553 ? _GEN_2703 : _GEN_2671; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2743 = _T_553 ? _GEN_2704 : _GEN_2672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2744 = _T_553 ? _GEN_2705 : _GEN_2673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2745 = _T_553 ? _GEN_2706 : _GEN_2674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2746 = _T_553 ? _GEN_2707 : _GEN_2675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2747 = _T_553 ? _GEN_2708 : _GEN_2676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2748 = _T_553 ? _GEN_2709 : _GEN_2677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2749 = _T_553 ? _GEN_2710 : _GEN_2678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2750 = _T_553 ? _GEN_2711 : _GEN_2679; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2751 = _T_553 ? _GEN_2712 : _GEN_2680; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2752 = _T_553 ? _GEN_2713 : _GEN_2681; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2753 = _T_553 ? _GEN_2714 : _GEN_2682; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2754 = _T_553 ? _GEN_2715 : _GEN_2683; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2755 = _T_553 ? _GEN_2716 : _GEN_2684; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2756 = _T_553 ? _GEN_2717 : _GEN_2685; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2757 = _T_553 ? _GEN_2718 : _GEN_2686; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2758 = _T_553 ? _GEN_2719 : _GEN_2687; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2759 = _T_553 ? _GEN_2720 : _GEN_2688; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2760 = _T_553 ? _GEN_2721 : _GEN_2689; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2761 = _T_553 ? _GEN_2722 : _GEN_2690; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [31:0] _GEN_2762 = _T_553 ? _GEN_2723 : _GEN_2691; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [6:0] _funct7_T_13 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_40 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_565 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_50 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_21 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _next_reg_T_94 = _GEN_31 * _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:65]
  wire [31:0] _next_reg_T_95 = _next_reg_T_80[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:80]
  wire [31:0] _next_reg_rd_30 = _next_reg_T_80[63:32]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:80]
  wire [31:0] _GEN_2763 = 5'h0 == rd ? _next_reg_T_80[63:32] : _GEN_2731; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2764 = 5'h1 == rd ? _next_reg_T_80[63:32] : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2765 = 5'h2 == rd ? _next_reg_T_80[63:32] : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2766 = 5'h3 == rd ? _next_reg_T_80[63:32] : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2767 = 5'h4 == rd ? _next_reg_T_80[63:32] : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2768 = 5'h5 == rd ? _next_reg_T_80[63:32] : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2769 = 5'h6 == rd ? _next_reg_T_80[63:32] : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2770 = 5'h7 == rd ? _next_reg_T_80[63:32] : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2771 = 5'h8 == rd ? _next_reg_T_80[63:32] : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2772 = 5'h9 == rd ? _next_reg_T_80[63:32] : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2773 = 5'ha == rd ? _next_reg_T_80[63:32] : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2774 = 5'hb == rd ? _next_reg_T_80[63:32] : _GEN_2742; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2775 = 5'hc == rd ? _next_reg_T_80[63:32] : _GEN_2743; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2776 = 5'hd == rd ? _next_reg_T_80[63:32] : _GEN_2744; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2777 = 5'he == rd ? _next_reg_T_80[63:32] : _GEN_2745; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2778 = 5'hf == rd ? _next_reg_T_80[63:32] : _GEN_2746; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2779 = 5'h10 == rd ? _next_reg_T_80[63:32] : _GEN_2747; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2780 = 5'h11 == rd ? _next_reg_T_80[63:32] : _GEN_2748; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2781 = 5'h12 == rd ? _next_reg_T_80[63:32] : _GEN_2749; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2782 = 5'h13 == rd ? _next_reg_T_80[63:32] : _GEN_2750; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2783 = 5'h14 == rd ? _next_reg_T_80[63:32] : _GEN_2751; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2784 = 5'h15 == rd ? _next_reg_T_80[63:32] : _GEN_2752; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2785 = 5'h16 == rd ? _next_reg_T_80[63:32] : _GEN_2753; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2786 = 5'h17 == rd ? _next_reg_T_80[63:32] : _GEN_2754; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2787 = 5'h18 == rd ? _next_reg_T_80[63:32] : _GEN_2755; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2788 = 5'h19 == rd ? _next_reg_T_80[63:32] : _GEN_2756; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2789 = 5'h1a == rd ? _next_reg_T_80[63:32] : _GEN_2757; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2790 = 5'h1b == rd ? _next_reg_T_80[63:32] : _GEN_2758; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2791 = 5'h1c == rd ? _next_reg_T_80[63:32] : _GEN_2759; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2792 = 5'h1d == rd ? _next_reg_T_80[63:32] : _GEN_2760; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2793 = 5'h1e == rd ? _next_reg_T_80[63:32] : _GEN_2761; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [31:0] _GEN_2794 = 5'h1f == rd ? _next_reg_T_80[63:32] : _GEN_2762; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [6:0] _GEN_2796 = _T_560 ? inst[31:25] : _GEN_2725; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2799 = _T_560 ? inst[14:12] : _GEN_2728; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2801 = _T_560 ? inst[6:0] : _GEN_2730; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2802 = _T_560 ? _GEN_2763 : _GEN_2731; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2803 = _T_560 ? _GEN_2764 : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2804 = _T_560 ? _GEN_2765 : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2805 = _T_560 ? _GEN_2766 : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2806 = _T_560 ? _GEN_2767 : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2807 = _T_560 ? _GEN_2768 : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2808 = _T_560 ? _GEN_2769 : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2809 = _T_560 ? _GEN_2770 : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2810 = _T_560 ? _GEN_2771 : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2811 = _T_560 ? _GEN_2772 : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2812 = _T_560 ? _GEN_2773 : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2813 = _T_560 ? _GEN_2774 : _GEN_2742; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2814 = _T_560 ? _GEN_2775 : _GEN_2743; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2815 = _T_560 ? _GEN_2776 : _GEN_2744; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2816 = _T_560 ? _GEN_2777 : _GEN_2745; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2817 = _T_560 ? _GEN_2778 : _GEN_2746; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2818 = _T_560 ? _GEN_2779 : _GEN_2747; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2819 = _T_560 ? _GEN_2780 : _GEN_2748; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2820 = _T_560 ? _GEN_2781 : _GEN_2749; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2821 = _T_560 ? _GEN_2782 : _GEN_2750; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2822 = _T_560 ? _GEN_2783 : _GEN_2751; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2823 = _T_560 ? _GEN_2784 : _GEN_2752; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2824 = _T_560 ? _GEN_2785 : _GEN_2753; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2825 = _T_560 ? _GEN_2786 : _GEN_2754; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2826 = _T_560 ? _GEN_2787 : _GEN_2755; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2827 = _T_560 ? _GEN_2788 : _GEN_2756; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2828 = _T_560 ? _GEN_2789 : _GEN_2757; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2829 = _T_560 ? _GEN_2790 : _GEN_2758; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2830 = _T_560 ? _GEN_2791 : _GEN_2759; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2831 = _T_560 ? _GEN_2792 : _GEN_2760; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2832 = _T_560 ? _GEN_2793 : _GEN_2761; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [31:0] _GEN_2833 = _T_560 ? _GEN_2794 : _GEN_2762; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [6:0] _funct7_T_14 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_41 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_572 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_51 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_96 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:16]
  wire [31:0] _now_reg_rs2_22 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_97 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:34]
  wire [32:0] _next_reg_T_98 = $signed(_T_300) / $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:23]
  wire [31:0] _next_reg_T_99 = _next_reg_T_98[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:41]
  wire [31:0] _now_reg_rs2_23 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_100 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:19]
  wire [31:0] _next_reg_T_101 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:99]
  wire [31:0] _next_reg_T_102 = 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:45]
  wire [32:0] _next_reg_T_103 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire [31:0] _next_reg_T_104 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire [31:0] _now_reg_rs1_52 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _next_reg_T_105 = _GEN_31 == _next_reg_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:18]
  wire [31:0] _next_reg_T_106 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:78]
  wire [31:0] _now_reg_rs2_24 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_107 = _GEN_840 == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:64]
  wire  _next_reg_T_108 = _GEN_31 == _next_reg_T_104 & _GEN_840 == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:52]
  wire [31:0] _next_reg_T_109 = 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:112]
  wire [32:0] _next_reg_T_110 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:89]
  wire [31:0] _next_reg_T_111 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:89]
  wire [31:0] _next_reg_T_112 = _next_reg_T_108 ? _next_reg_T_104 : _next_reg_T_98[31:0]; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_T_113 = _next_reg_T_100 ? 32'hffffffff : _next_reg_T_112; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_31 = _next_reg_T_100 ? 32'hffffffff : _next_reg_T_112; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_2834 = 5'h0 == rd ? _next_reg_T_113 : _GEN_2802; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2835 = 5'h1 == rd ? _next_reg_T_113 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2836 = 5'h2 == rd ? _next_reg_T_113 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2837 = 5'h3 == rd ? _next_reg_T_113 : _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2838 = 5'h4 == rd ? _next_reg_T_113 : _GEN_2806; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2839 = 5'h5 == rd ? _next_reg_T_113 : _GEN_2807; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2840 = 5'h6 == rd ? _next_reg_T_113 : _GEN_2808; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2841 = 5'h7 == rd ? _next_reg_T_113 : _GEN_2809; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2842 = 5'h8 == rd ? _next_reg_T_113 : _GEN_2810; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2843 = 5'h9 == rd ? _next_reg_T_113 : _GEN_2811; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2844 = 5'ha == rd ? _next_reg_T_113 : _GEN_2812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2845 = 5'hb == rd ? _next_reg_T_113 : _GEN_2813; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2846 = 5'hc == rd ? _next_reg_T_113 : _GEN_2814; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2847 = 5'hd == rd ? _next_reg_T_113 : _GEN_2815; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2848 = 5'he == rd ? _next_reg_T_113 : _GEN_2816; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2849 = 5'hf == rd ? _next_reg_T_113 : _GEN_2817; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2850 = 5'h10 == rd ? _next_reg_T_113 : _GEN_2818; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2851 = 5'h11 == rd ? _next_reg_T_113 : _GEN_2819; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2852 = 5'h12 == rd ? _next_reg_T_113 : _GEN_2820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2853 = 5'h13 == rd ? _next_reg_T_113 : _GEN_2821; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2854 = 5'h14 == rd ? _next_reg_T_113 : _GEN_2822; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2855 = 5'h15 == rd ? _next_reg_T_113 : _GEN_2823; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2856 = 5'h16 == rd ? _next_reg_T_113 : _GEN_2824; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2857 = 5'h17 == rd ? _next_reg_T_113 : _GEN_2825; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2858 = 5'h18 == rd ? _next_reg_T_113 : _GEN_2826; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2859 = 5'h19 == rd ? _next_reg_T_113 : _GEN_2827; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2860 = 5'h1a == rd ? _next_reg_T_113 : _GEN_2828; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2861 = 5'h1b == rd ? _next_reg_T_113 : _GEN_2829; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2862 = 5'h1c == rd ? _next_reg_T_113 : _GEN_2830; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2863 = 5'h1d == rd ? _next_reg_T_113 : _GEN_2831; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2864 = 5'h1e == rd ? _next_reg_T_113 : _GEN_2832; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [31:0] _GEN_2865 = 5'h1f == rd ? _next_reg_T_113 : _GEN_2833; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [6:0] _GEN_2867 = _T_567 ? inst[31:25] : _GEN_2796; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2870 = _T_567 ? inst[14:12] : _GEN_2799; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2872 = _T_567 ? inst[6:0] : _GEN_2801; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2873 = _T_567 ? _GEN_2834 : _GEN_2802; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2874 = _T_567 ? _GEN_2835 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2875 = _T_567 ? _GEN_2836 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2876 = _T_567 ? _GEN_2837 : _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2877 = _T_567 ? _GEN_2838 : _GEN_2806; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2878 = _T_567 ? _GEN_2839 : _GEN_2807; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2879 = _T_567 ? _GEN_2840 : _GEN_2808; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2880 = _T_567 ? _GEN_2841 : _GEN_2809; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2881 = _T_567 ? _GEN_2842 : _GEN_2810; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2882 = _T_567 ? _GEN_2843 : _GEN_2811; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2883 = _T_567 ? _GEN_2844 : _GEN_2812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2884 = _T_567 ? _GEN_2845 : _GEN_2813; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2885 = _T_567 ? _GEN_2846 : _GEN_2814; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2886 = _T_567 ? _GEN_2847 : _GEN_2815; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2887 = _T_567 ? _GEN_2848 : _GEN_2816; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2888 = _T_567 ? _GEN_2849 : _GEN_2817; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2889 = _T_567 ? _GEN_2850 : _GEN_2818; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2890 = _T_567 ? _GEN_2851 : _GEN_2819; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2891 = _T_567 ? _GEN_2852 : _GEN_2820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2892 = _T_567 ? _GEN_2853 : _GEN_2821; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2893 = _T_567 ? _GEN_2854 : _GEN_2822; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2894 = _T_567 ? _GEN_2855 : _GEN_2823; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2895 = _T_567 ? _GEN_2856 : _GEN_2824; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2896 = _T_567 ? _GEN_2857 : _GEN_2825; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2897 = _T_567 ? _GEN_2858 : _GEN_2826; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2898 = _T_567 ? _GEN_2859 : _GEN_2827; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2899 = _T_567 ? _GEN_2860 : _GEN_2828; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2900 = _T_567 ? _GEN_2861 : _GEN_2829; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2901 = _T_567 ? _GEN_2862 : _GEN_2830; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2902 = _T_567 ? _GEN_2863 : _GEN_2831; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2903 = _T_567 ? _GEN_2864 : _GEN_2832; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [31:0] _GEN_2904 = _T_567 ? _GEN_2865 : _GEN_2833; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [6:0] _funct7_T_15 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_42 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_579 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_53 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_25 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_114 = _GEN_31 / _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 58:15]
  wire [31:0] _now_reg_rs2_26 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_115 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 60:19]
  wire [31:0] _next_reg_T_116 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 60:40]
  wire [31:0] _next_reg_T_117 = _next_reg_T_100 ? 32'hffffffff : _next_reg_T_114; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_32 = _next_reg_T_100 ? 32'hffffffff : _next_reg_T_114; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_2905 = 5'h0 == rd ? _next_reg_T_117 : _GEN_2873; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2906 = 5'h1 == rd ? _next_reg_T_117 : _GEN_2874; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2907 = 5'h2 == rd ? _next_reg_T_117 : _GEN_2875; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2908 = 5'h3 == rd ? _next_reg_T_117 : _GEN_2876; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2909 = 5'h4 == rd ? _next_reg_T_117 : _GEN_2877; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2910 = 5'h5 == rd ? _next_reg_T_117 : _GEN_2878; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2911 = 5'h6 == rd ? _next_reg_T_117 : _GEN_2879; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2912 = 5'h7 == rd ? _next_reg_T_117 : _GEN_2880; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2913 = 5'h8 == rd ? _next_reg_T_117 : _GEN_2881; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2914 = 5'h9 == rd ? _next_reg_T_117 : _GEN_2882; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2915 = 5'ha == rd ? _next_reg_T_117 : _GEN_2883; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2916 = 5'hb == rd ? _next_reg_T_117 : _GEN_2884; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2917 = 5'hc == rd ? _next_reg_T_117 : _GEN_2885; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2918 = 5'hd == rd ? _next_reg_T_117 : _GEN_2886; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2919 = 5'he == rd ? _next_reg_T_117 : _GEN_2887; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2920 = 5'hf == rd ? _next_reg_T_117 : _GEN_2888; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2921 = 5'h10 == rd ? _next_reg_T_117 : _GEN_2889; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2922 = 5'h11 == rd ? _next_reg_T_117 : _GEN_2890; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2923 = 5'h12 == rd ? _next_reg_T_117 : _GEN_2891; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2924 = 5'h13 == rd ? _next_reg_T_117 : _GEN_2892; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2925 = 5'h14 == rd ? _next_reg_T_117 : _GEN_2893; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2926 = 5'h15 == rd ? _next_reg_T_117 : _GEN_2894; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2927 = 5'h16 == rd ? _next_reg_T_117 : _GEN_2895; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2928 = 5'h17 == rd ? _next_reg_T_117 : _GEN_2896; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2929 = 5'h18 == rd ? _next_reg_T_117 : _GEN_2897; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2930 = 5'h19 == rd ? _next_reg_T_117 : _GEN_2898; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2931 = 5'h1a == rd ? _next_reg_T_117 : _GEN_2899; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2932 = 5'h1b == rd ? _next_reg_T_117 : _GEN_2900; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2933 = 5'h1c == rd ? _next_reg_T_117 : _GEN_2901; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2934 = 5'h1d == rd ? _next_reg_T_117 : _GEN_2902; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2935 = 5'h1e == rd ? _next_reg_T_117 : _GEN_2903; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [31:0] _GEN_2936 = 5'h1f == rd ? _next_reg_T_117 : _GEN_2904; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [6:0] _GEN_2938 = _T_574 ? inst[31:25] : _GEN_2867; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_2941 = _T_574 ? inst[14:12] : _GEN_2870; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2943 = _T_574 ? inst[6:0] : _GEN_2872; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_2944 = _T_574 ? _GEN_2905 : _GEN_2873; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2945 = _T_574 ? _GEN_2906 : _GEN_2874; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2946 = _T_574 ? _GEN_2907 : _GEN_2875; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2947 = _T_574 ? _GEN_2908 : _GEN_2876; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2948 = _T_574 ? _GEN_2909 : _GEN_2877; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2949 = _T_574 ? _GEN_2910 : _GEN_2878; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2950 = _T_574 ? _GEN_2911 : _GEN_2879; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2951 = _T_574 ? _GEN_2912 : _GEN_2880; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2952 = _T_574 ? _GEN_2913 : _GEN_2881; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2953 = _T_574 ? _GEN_2914 : _GEN_2882; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2954 = _T_574 ? _GEN_2915 : _GEN_2883; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2955 = _T_574 ? _GEN_2916 : _GEN_2884; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2956 = _T_574 ? _GEN_2917 : _GEN_2885; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2957 = _T_574 ? _GEN_2918 : _GEN_2886; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2958 = _T_574 ? _GEN_2919 : _GEN_2887; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2959 = _T_574 ? _GEN_2920 : _GEN_2888; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2960 = _T_574 ? _GEN_2921 : _GEN_2889; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2961 = _T_574 ? _GEN_2922 : _GEN_2890; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2962 = _T_574 ? _GEN_2923 : _GEN_2891; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2963 = _T_574 ? _GEN_2924 : _GEN_2892; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2964 = _T_574 ? _GEN_2925 : _GEN_2893; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2965 = _T_574 ? _GEN_2926 : _GEN_2894; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2966 = _T_574 ? _GEN_2927 : _GEN_2895; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2967 = _T_574 ? _GEN_2928 : _GEN_2896; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2968 = _T_574 ? _GEN_2929 : _GEN_2897; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2969 = _T_574 ? _GEN_2930 : _GEN_2898; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2970 = _T_574 ? _GEN_2931 : _GEN_2899; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2971 = _T_574 ? _GEN_2932 : _GEN_2900; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2972 = _T_574 ? _GEN_2933 : _GEN_2901; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2973 = _T_574 ? _GEN_2934 : _GEN_2902; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2974 = _T_574 ? _GEN_2935 : _GEN_2903; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [31:0] _GEN_2975 = _T_574 ? _GEN_2936 : _GEN_2904; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [6:0] _funct7_T_16 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_43 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_586 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_54 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_118 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:16]
  wire [31:0] _now_reg_rs2_27 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_119 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:34]
  wire [31:0] _next_reg_T_120 = $signed(_T_300) % $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:23]
  wire [31:0] _next_reg_T_121 = $signed(_T_300) % $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:42]
  wire [31:0] _now_reg_rs2_28 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_122 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 68:19]
  wire [31:0] _next_reg_T_123 = 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:45]
  wire [32:0] _next_reg_T_124 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:22]
  wire [31:0] _next_reg_T_125 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:22]
  wire [31:0] _now_reg_rs1_55 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire  _next_reg_T_126 = _GEN_31 == _next_reg_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:18]
  wire [31:0] _next_reg_T_127 = 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:78]
  wire [31:0] _now_reg_rs2_29 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_128 = _GEN_840 == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:64]
  wire  _next_reg_T_129 = _next_reg_T_105 & _next_reg_T_107; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 69:52]
  wire [31:0] _next_reg_T_130 = _next_reg_T_108 ? 32'h0 : _next_reg_T_121; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _now_reg_rs1_56 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_131 = _next_reg_T_100 ? _GEN_31 : _next_reg_T_130; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_33 = _next_reg_T_100 ? _GEN_31 : _next_reg_T_130; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_2976 = 5'h0 == rd ? _next_reg_T_131 : _GEN_2944; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2977 = 5'h1 == rd ? _next_reg_T_131 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2978 = 5'h2 == rd ? _next_reg_T_131 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2979 = 5'h3 == rd ? _next_reg_T_131 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2980 = 5'h4 == rd ? _next_reg_T_131 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2981 = 5'h5 == rd ? _next_reg_T_131 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2982 = 5'h6 == rd ? _next_reg_T_131 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2983 = 5'h7 == rd ? _next_reg_T_131 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2984 = 5'h8 == rd ? _next_reg_T_131 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2985 = 5'h9 == rd ? _next_reg_T_131 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2986 = 5'ha == rd ? _next_reg_T_131 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2987 = 5'hb == rd ? _next_reg_T_131 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2988 = 5'hc == rd ? _next_reg_T_131 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2989 = 5'hd == rd ? _next_reg_T_131 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2990 = 5'he == rd ? _next_reg_T_131 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2991 = 5'hf == rd ? _next_reg_T_131 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2992 = 5'h10 == rd ? _next_reg_T_131 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2993 = 5'h11 == rd ? _next_reg_T_131 : _GEN_2961; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2994 = 5'h12 == rd ? _next_reg_T_131 : _GEN_2962; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2995 = 5'h13 == rd ? _next_reg_T_131 : _GEN_2963; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2996 = 5'h14 == rd ? _next_reg_T_131 : _GEN_2964; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2997 = 5'h15 == rd ? _next_reg_T_131 : _GEN_2965; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2998 = 5'h16 == rd ? _next_reg_T_131 : _GEN_2966; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_2999 = 5'h17 == rd ? _next_reg_T_131 : _GEN_2967; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3000 = 5'h18 == rd ? _next_reg_T_131 : _GEN_2968; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3001 = 5'h19 == rd ? _next_reg_T_131 : _GEN_2969; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3002 = 5'h1a == rd ? _next_reg_T_131 : _GEN_2970; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3003 = 5'h1b == rd ? _next_reg_T_131 : _GEN_2971; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3004 = 5'h1c == rd ? _next_reg_T_131 : _GEN_2972; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3005 = 5'h1d == rd ? _next_reg_T_131 : _GEN_2973; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3006 = 5'h1e == rd ? _next_reg_T_131 : _GEN_2974; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [31:0] _GEN_3007 = 5'h1f == rd ? _next_reg_T_131 : _GEN_2975; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [6:0] _GEN_3009 = _T_581 ? inst[31:25] : _GEN_2938; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3012 = _T_581 ? inst[14:12] : _GEN_2941; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3014 = _T_581 ? inst[6:0] : _GEN_2943; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3015 = _T_581 ? _GEN_2976 : _GEN_2944; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3016 = _T_581 ? _GEN_2977 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3017 = _T_581 ? _GEN_2978 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3018 = _T_581 ? _GEN_2979 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3019 = _T_581 ? _GEN_2980 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3020 = _T_581 ? _GEN_2981 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3021 = _T_581 ? _GEN_2982 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3022 = _T_581 ? _GEN_2983 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3023 = _T_581 ? _GEN_2984 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3024 = _T_581 ? _GEN_2985 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3025 = _T_581 ? _GEN_2986 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3026 = _T_581 ? _GEN_2987 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3027 = _T_581 ? _GEN_2988 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3028 = _T_581 ? _GEN_2989 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3029 = _T_581 ? _GEN_2990 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3030 = _T_581 ? _GEN_2991 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3031 = _T_581 ? _GEN_2992 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3032 = _T_581 ? _GEN_2993 : _GEN_2961; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3033 = _T_581 ? _GEN_2994 : _GEN_2962; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3034 = _T_581 ? _GEN_2995 : _GEN_2963; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3035 = _T_581 ? _GEN_2996 : _GEN_2964; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3036 = _T_581 ? _GEN_2997 : _GEN_2965; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3037 = _T_581 ? _GEN_2998 : _GEN_2966; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3038 = _T_581 ? _GEN_2999 : _GEN_2967; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3039 = _T_581 ? _GEN_3000 : _GEN_2968; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3040 = _T_581 ? _GEN_3001 : _GEN_2969; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3041 = _T_581 ? _GEN_3002 : _GEN_2970; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3042 = _T_581 ? _GEN_3003 : _GEN_2971; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3043 = _T_581 ? _GEN_3004 : _GEN_2972; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3044 = _T_581 ? _GEN_3005 : _GEN_2973; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3045 = _T_581 ? _GEN_3006 : _GEN_2974; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [31:0] _GEN_3046 = _T_581 ? _GEN_3007 : _GEN_2975; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [6:0] _funct7_T_17 = inst[31:25]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [2:0] _funct3_T_44 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_593 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _now_reg_rs1_57 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _now_reg_rs2_30 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [31:0] _next_reg_T_132 = _GEN_31 % _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 75:15]
  wire [31:0] _now_reg_rs2_31 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire  _next_reg_T_133 = _GEN_840 == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 77:19]
  wire [31:0] _now_reg_rs1_58 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [31:0] _next_reg_T_134 = _next_reg_T_100 ? _GEN_31 : _next_reg_T_132; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_rd_34 = _next_reg_T_100 ? _GEN_31 : _next_reg_T_132; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _GEN_3047 = 5'h0 == rd ? _next_reg_T_134 : _GEN_3015; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3048 = 5'h1 == rd ? _next_reg_T_134 : _GEN_3016; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3049 = 5'h2 == rd ? _next_reg_T_134 : _GEN_3017; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3050 = 5'h3 == rd ? _next_reg_T_134 : _GEN_3018; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3051 = 5'h4 == rd ? _next_reg_T_134 : _GEN_3019; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3052 = 5'h5 == rd ? _next_reg_T_134 : _GEN_3020; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3053 = 5'h6 == rd ? _next_reg_T_134 : _GEN_3021; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3054 = 5'h7 == rd ? _next_reg_T_134 : _GEN_3022; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3055 = 5'h8 == rd ? _next_reg_T_134 : _GEN_3023; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3056 = 5'h9 == rd ? _next_reg_T_134 : _GEN_3024; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3057 = 5'ha == rd ? _next_reg_T_134 : _GEN_3025; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3058 = 5'hb == rd ? _next_reg_T_134 : _GEN_3026; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3059 = 5'hc == rd ? _next_reg_T_134 : _GEN_3027; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3060 = 5'hd == rd ? _next_reg_T_134 : _GEN_3028; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3061 = 5'he == rd ? _next_reg_T_134 : _GEN_3029; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3062 = 5'hf == rd ? _next_reg_T_134 : _GEN_3030; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3063 = 5'h10 == rd ? _next_reg_T_134 : _GEN_3031; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3064 = 5'h11 == rd ? _next_reg_T_134 : _GEN_3032; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3065 = 5'h12 == rd ? _next_reg_T_134 : _GEN_3033; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3066 = 5'h13 == rd ? _next_reg_T_134 : _GEN_3034; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3067 = 5'h14 == rd ? _next_reg_T_134 : _GEN_3035; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3068 = 5'h15 == rd ? _next_reg_T_134 : _GEN_3036; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3069 = 5'h16 == rd ? _next_reg_T_134 : _GEN_3037; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3070 = 5'h17 == rd ? _next_reg_T_134 : _GEN_3038; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3071 = 5'h18 == rd ? _next_reg_T_134 : _GEN_3039; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3072 = 5'h19 == rd ? _next_reg_T_134 : _GEN_3040; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3073 = 5'h1a == rd ? _next_reg_T_134 : _GEN_3041; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3074 = 5'h1b == rd ? _next_reg_T_134 : _GEN_3042; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3075 = 5'h1c == rd ? _next_reg_T_134 : _GEN_3043; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3076 = 5'h1d == rd ? _next_reg_T_134 : _GEN_3044; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3077 = 5'h1e == rd ? _next_reg_T_134 : _GEN_3045; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [31:0] _GEN_3078 = 5'h1f == rd ? _next_reg_T_134 : _GEN_3046; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [6:0] _GEN_3080 = _T_588 ? inst[31:25] : _GEN_3009; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_3083 = _T_588 ? inst[14:12] : _GEN_3012; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3085 = _T_588 ? inst[6:0] : _GEN_3014; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] _GEN_3086 = _T_588 ? _GEN_3047 : _GEN_3015; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3087 = _T_588 ? _GEN_3048 : _GEN_3016; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3088 = _T_588 ? _GEN_3049 : _GEN_3017; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3089 = _T_588 ? _GEN_3050 : _GEN_3018; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3090 = _T_588 ? _GEN_3051 : _GEN_3019; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3091 = _T_588 ? _GEN_3052 : _GEN_3020; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3092 = _T_588 ? _GEN_3053 : _GEN_3021; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3093 = _T_588 ? _GEN_3054 : _GEN_3022; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3094 = _T_588 ? _GEN_3055 : _GEN_3023; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3095 = _T_588 ? _GEN_3056 : _GEN_3024; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3096 = _T_588 ? _GEN_3057 : _GEN_3025; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3097 = _T_588 ? _GEN_3058 : _GEN_3026; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3098 = _T_588 ? _GEN_3059 : _GEN_3027; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3099 = _T_588 ? _GEN_3060 : _GEN_3028; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3100 = _T_588 ? _GEN_3061 : _GEN_3029; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3101 = _T_588 ? _GEN_3062 : _GEN_3030; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3102 = _T_588 ? _GEN_3063 : _GEN_3031; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3103 = _T_588 ? _GEN_3064 : _GEN_3032; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3104 = _T_588 ? _GEN_3065 : _GEN_3033; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3105 = _T_588 ? _GEN_3066 : _GEN_3034; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3106 = _T_588 ? _GEN_3067 : _GEN_3035; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3107 = _T_588 ? _GEN_3068 : _GEN_3036; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3108 = _T_588 ? _GEN_3069 : _GEN_3037; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3109 = _T_588 ? _GEN_3070 : _GEN_3038; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3110 = _T_588 ? _GEN_3071 : _GEN_3039; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3111 = _T_588 ? _GEN_3072 : _GEN_3040; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3112 = _T_588 ? _GEN_3073 : _GEN_3041; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3113 = _T_588 ? _GEN_3074 : _GEN_3042; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3114 = _T_588 ? _GEN_3075 : _GEN_3043; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3115 = _T_588 ? _GEN_3076 : _GEN_3044; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3116 = _T_588 ? _GEN_3077 : _GEN_3045; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [31:0] _GEN_3117 = _T_588 ? _GEN_3078 : _GEN_3046; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [2:0] _funct3_T_45 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_599 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire  mstatusOld_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [7:0] mstatusOld_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [31:0] _mstatusNew_WIRE_1 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusNew_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_1 = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_5 = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_8 = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] mstatusNew_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_13 = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [7:0] mstatusNew_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusOld_WIRE_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_8 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _next_internal_privilegeMode_T = {1'h0,mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 125:41]
  wire  _mstatusNew_WIRE_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusOld_WIRE_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_5 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusNew_sie = illegalSret | illegalSModeSret ? mstatusOld_sie : mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 124:35]
  wire  _GEN_3120 = mstatusNew_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 124:35]
  wire  _mstatusNew_WIRE_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] next_csr_mstatus_lo_lo_lo = {mstatusNew_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_4 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_3 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi = {mstatusOld_pad2,mstatusOld_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_2 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [2:0] next_csr_mstatus_lo_lo_hi = {mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [4:0] next_csr_mstatus_lo_lo = {mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3,mstatusNew_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_6 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_spie = illegalSret | illegalSModeSret ? mstatusOld_spie : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 126:35]
  wire  _GEN_3122 = mstatusNew_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 126:35]
  wire [1:0] next_csr_mstatus_lo_hi_lo = {mstatusOld_ube,mstatusNew_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [1:0] _mstatusNew_WIRE_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_9 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_spp = (illegalSret | illegalSModeSret) & mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 127:35]
  wire  _GEN_3123 = mstatusNew_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 127:35]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi = {mstatusOld_vs,mstatusNew_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_7 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [3:0] next_csr_mstatus_lo_hi_hi = {mstatusOld_vs,mstatusNew_spp,mstatusOld_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [5:0] next_csr_mstatus_lo_hi = {mstatusOld_vs,mstatusNew_spp,mstatusOld_mpie,mstatusOld_ube,mstatusNew_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [10:0] next_csr_mstatus_lo = {mstatusOld_vs,mstatusNew_spp,mstatusOld_mpie,mstatusOld_ube,mstatusNew_spie,
    mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3,mstatusNew_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [1:0] _mstatusNew_WIRE_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_11 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_WIRE_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_10 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [3:0] next_csr_mstatus_hi_lo_lo = {mstatusOld_fs,mstatusOld_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_14 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  mstatusNew_mprv = (illegalSret | illegalSModeSret) & mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 128:35]
  wire  _GEN_3124 = mstatusNew_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 128:35]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi = {mstatusOld_sum,mstatusNew_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [1:0] _mstatusNew_WIRE_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] _mstatusNew_T_12 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [3:0] next_csr_mstatus_hi_lo_hi = {mstatusOld_sum,mstatusNew_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [7:0] next_csr_mstatus_hi_lo = {mstatusOld_sum,mstatusNew_mprv,mstatusOld_xs,mstatusOld_fs,mstatusOld_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_17 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_WIRE_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_16 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_15 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [2:0] next_csr_mstatus_hi_hi_lo = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_20 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [7:0] _mstatusNew_WIRE_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [7:0] _mstatusNew_T_19 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _mstatusNew_WIRE_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire  _mstatusNew_T_18 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:55]
  wire [9:0] next_csr_mstatus_hi_hi_hi = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [12:0] next_csr_mstatus_hi_hi = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [20:0] next_csr_mstatus_hi = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [31:0] _next_csr_mstatus_T = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo,next_csr_mstatus_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _GEN_3119 = illegalSret | illegalSModeSret | _GEN_2540; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3137 = _T_595 ? _GEN_3119 : _GEN_2540; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire  _GEN_3149 = io_now_internal_privilegeMode == 2'h3 ? _GEN_3137 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3163 = _T_602 ? _GEN_3149 : _GEN_3137; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_3180 = illegalInstruction | _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 145:33]
  wire  raiseExceptionIntr = io_valid & _GEN_3180; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire  _GEN_3308 = raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [31:0] now_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _delegS_T = io_now_csr_medeleg >> exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:24]
  wire  _delegS_T_1 = _delegS_T[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:24]
  wire  _delegS_T_2 = io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:70]
  wire  delegS = _delegS_T[0] & io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:39]
  wire [7:0] now_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_621 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] now_csr_sepc = io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3195 = 8'h20 == io_now_csr_MXLEN ? io_now_pc : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 254:35]
  wire [31:0] _GEN_3230 = delegS ? _GEN_3195 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_3247 = raiseExceptionIntr ? _GEN_3230 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_sepc = io_valid ? _GEN_3247 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3336 = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _retTarget_T = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [1:0] _GEN_3121 = illegalSret | illegalSModeSret ? io_now_internal_privilegeMode : _next_internal_privilegeMode_T
    ; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 125:35]
  wire [31:0] _GEN_3125 = illegalSret | illegalSModeSret ? io_now_csr_mstatus : _next_csr_mstatus_T; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 129:35]
  wire [31:0] _GEN_3126 = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  _GEN_3127 = illegalSret | illegalSModeSret ? _GEN_1923 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 132:25]
  wire [31:0] _GEN_3128 = illegalSret | illegalSModeSret ? _GEN_1924 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 133:25]
  wire [2:0] _GEN_3132 = _T_595 ? inst[14:12] : _GEN_3083; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3134 = _T_595 ? inst[6:0] : _GEN_3085; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [1:0] _GEN_3138 = _T_595 ? _GEN_3121 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_3139 = _T_595 ? _GEN_3125 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_3140 = next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  _GEN_3141 = _T_595 ? _GEN_3127 : _GEN_1923; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [31:0] _GEN_3142 = _T_595 ? _GEN_3128 : _GEN_1924; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [2:0] _funct3_T_46 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_606 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [31:0] _mstatusOld_WIRE_3 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusOld_1_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] mstatusOld_1_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [7:0] mstatusOld_1_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusOld_1_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [31:0] _mstatusNew_WIRE_3 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusNew_1_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_24 = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_28 = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_31 = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [7:0] mstatusNew_1_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  mstatusNew_1_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_22 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_21 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_lo_lo_lo_1 = {mstatusOld_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_25 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusOld_WIRE_2_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_28 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  mstatusNew_1_mie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_1 = {mstatusOld_pad2,mstatusOld_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_23 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [2:0] next_csr_mstatus_lo_lo_hi_1 = {mstatusOld_pad2,mstatusOld_mpie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [4:0] next_csr_mstatus_lo_lo_1 = {mstatusOld_pad2,mstatusOld_mpie,mstatusOld_pad3,mstatusOld_sie,mstatusOld_pad4}
    ; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_27 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_26 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_lo_hi_lo_1 = {mstatusOld_ube,mstatusOld_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [1:0] _mstatusNew_WIRE_2_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_30 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_29 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_1 = {mstatusOld_vs,mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  mstatusNew_1_mpie = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:32 93:35]
  wire [3:0] next_csr_mstatus_lo_hi_hi_1 = {mstatusOld_vs,mstatusOld_spp,1'h1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [5:0] next_csr_mstatus_lo_hi_1 = {mstatusOld_vs,mstatusOld_spp,1'h1,mstatusOld_ube,mstatusOld_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [10:0] next_csr_mstatus_lo_1 = {mstatusOld_vs,mstatusOld_spp,1'h1,mstatusOld_ube,mstatusOld_spie,mstatusOld_pad2,
    mstatusOld_mpie,mstatusOld_pad3,mstatusOld_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [1:0] _mstatusNew_WIRE_2_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_32 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] mstatusNew_1_mpp = 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:32 98:24]
  wire [3:0] next_csr_mstatus_hi_lo_lo_1 = {mstatusOld_fs,2'h3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_35 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_34 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_1 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [1:0] _mstatusNew_WIRE_2_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] _mstatusNew_T_33 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [3:0] next_csr_mstatus_hi_lo_hi_1 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [7:0] next_csr_mstatus_hi_lo_1 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,2'h3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_38 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_37 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_1 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_36 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [2:0] next_csr_mstatus_hi_hi_lo_1 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_41 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [7:0] _mstatusNew_WIRE_2_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [7:0] _mstatusNew_T_40 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_1 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire  _mstatusNew_WIRE_2_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_T_39 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire [9:0] next_csr_mstatus_hi_hi_hi_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [12:0] next_csr_mstatus_hi_hi_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [20:0] next_csr_mstatus_hi_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [31:0] _next_csr_mstatus_T_1 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_1,next_csr_mstatus_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [31:0] now_csr_mepc = io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  _T_639 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_3215 = _T_621 ? io_now_pc : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 186:35]
  wire [31:0] _GEN_3239 = delegS ? io_now_csr_mepc : _GEN_3215; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_3253 = raiseExceptionIntr ? _GEN_3239 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_mepc = io_valid ? _GEN_3253 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3339 = next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _retTarget_T_1 = next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [1:0] _mstatusOld_WIRE_2_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_31 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _GEN_3143 = io_now_internal_privilegeMode == 2'h3 ? mstatusOld_mpp : _GEN_3138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 92:35]
  wire [31:0] _GEN_3144 = io_now_internal_privilegeMode == 2'h3 ? _next_csr_mstatus_T_1 : _GEN_3139; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:24 88:48]
  wire [31:0] _GEN_3145 = io_now_internal_privilegeMode == 2'h3 ? next_csr_mepc : next_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 101:24 88:48]
  wire  _GEN_3146 = io_now_internal_privilegeMode == 2'h3 | _GEN_3141; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 103:25 88:48]
  wire [31:0] _GEN_3147 = io_now_internal_privilegeMode == 2'h3 ? io_now_csr_mepc : _GEN_3142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 104:25 88:48]
  wire [2:0] _GEN_3153 = _T_602 ? inst[14:12] : _GEN_3132; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3155 = _T_602 ? inst[6:0] : _GEN_3134; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [1:0] _GEN_3157 = _T_602 ? _GEN_3143 : _GEN_3138; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _GEN_3158 = _T_602 ? _GEN_3144 : _GEN_3139; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] retTarget = _T_602 ? _GEN_3145 : next_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_3160 = _T_602 ? _GEN_3146 : _GEN_3141; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _GEN_3161 = _T_602 ? _GEN_3147 : _GEN_3142; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [2:0] _funct3_T_47 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_613 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_3167 = _T_609 ? inst[14:12] : _GEN_3153; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3169 = _T_609 ? inst[6:0] : _GEN_3155; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [2:0] _funct3_T_48 = inst[14:12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 31:23]
  wire [6:0] _T_619 = inst[6:0]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 32:33]
  wire [2:0] _GEN_3174 = _T_615 ? inst[14:12] : _GEN_3167; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3176 = _T_615 ? inst[6:0] : _GEN_3169; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 35:16]
  wire [31:0] now_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [1:0] _T_635 = io_now_csr_stvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:27]
  wire  _T_636 = 2'h0 == io_now_csr_stvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35]
  wire  _T_637 = 2'h1 == io_now_csr_stvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35]
  wire  _GEN_3190 = 2'h1 == io_now_csr_stvec[1:0] | _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 316:29]
  wire  _GEN_3192 = 2'h0 == io_now_csr_stvec[1:0] | _GEN_3190; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 311:29]
  wire  _GEN_3202 = 8'h20 == io_now_csr_MXLEN ? _GEN_3192 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] now_csr_mtvec = io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [1:0] _T_651 = io_now_csr_mtvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:27]
  wire  _T_652 = 2'h0 == io_now_csr_mtvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35]
  wire  _T_653 = 2'h1 == io_now_csr_mtvec[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35]
  wire  _GEN_3210 = 2'h1 == io_now_csr_mtvec[1:0] | _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 242:29]
  wire  _GEN_3212 = 2'h0 == io_now_csr_mtvec[1:0] | _GEN_3210; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 237:29]
  wire  _GEN_3222 = _T_621 ? _GEN_3212 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire  _GEN_3233 = delegS ? _GEN_3202 : _GEN_3222; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire  _GEN_3250 = raiseExceptionIntr ? _GEN_3233 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire  global_data_setpc = io_valid & _GEN_3250; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 113:21]
  wire  _GEN_3304 = global_data_setpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 113:21]
  wire  _T_620 = ~global_data_setpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 150:10]
  wire [32:0] _next_pc_T_18 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 156:27]
  wire [31:0] _next_pc_T_19 = io_now_pc + 32'h4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 156:27]
  wire [31:0] _GEN_3178 = ~global_data_setpc ? _next_reg_T_43 : _GEN_3161; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 150:30 156:17]
  wire [31:0] _event_exceptionInst_T = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _mstatusOld_WIRE_5 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusOld_2_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] mstatusOld_2_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [7:0] mstatusOld_2_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusOld_2_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [31:0] _mstatusNew_WIRE_5 = io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire  mstatusNew_2_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_43 = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_45 = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_47 = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_49 = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_50 = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] mstatusNew_2_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_52 = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] mstatusNew_2_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] mstatusNew_2_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [7:0] mstatusNew_2_pad0 = io_now_csr_mstatus[30:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_sd = io_now_csr_mstatus[31]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [30:0] _next_csr_scause_T = {26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_scause_T_1 = {1'h0,26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 252:29]
  wire  _GEN_3198 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 164:35 257:35]
  wire  _mstatusNew_WIRE_4_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_sie = delegS ? 1'h0 : mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_3227 = mstatusNew_2_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _mstatusNew_WIRE_4_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_42 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] next_csr_mstatus_lo_lo_lo_2 = {mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_46 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_WIRE_4_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _GEN_3218 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 174:35 189:35]
  wire  mstatusNew_2_mie = delegS & mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_3237 = mstatusNew_2_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_2 = {mstatusOld_pad2,mstatusNew_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_44 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [2:0] next_csr_mstatus_lo_lo_hi_2 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [4:0] next_csr_mstatus_lo_lo_2 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_48 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusOld_WIRE_4_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_43 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _GEN_3197 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusNew_WIRE_4_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  mstatusNew_2_spie = delegS ? mstatusOld_sie : mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_3226 = mstatusNew_2_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] next_csr_mstatus_lo_hi_lo_2 = {mstatusOld_ube,mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _mstatusNew_WIRE_4_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_51 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _GEN_3196 = io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 162:35 255:35]
  wire  _mstatusNew_WIRE_4_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _GEN_3225 = delegS ? io_now_internal_privilegeMode : {{1'd0}, mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_spp = _GEN_3225[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:30]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_2 = {mstatusOld_vs,mstatusNew_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusOld_WIRE_4_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_45 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _GEN_3217 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  mstatusNew_2_mpie = delegS ? mstatusOld_mpie : mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  _GEN_3236 = mstatusNew_2_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [3:0] next_csr_mstatus_lo_hi_hi_2 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [5:0] next_csr_mstatus_lo_hi_2 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,
    mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [10:0] next_csr_mstatus_lo_2 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,mstatusNew_2_spie
    ,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _mstatusNew_WIRE_4_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_53 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_WIRE_4_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _GEN_3216 = io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 172:35 187:35]
  wire [1:0] mstatusNew_2_mpp = delegS ? mstatusOld_mpp : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] _GEN_3235 = mstatusNew_2_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [3:0] next_csr_mstatus_hi_lo_lo_2 = {mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_56 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_WIRE_4_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_55 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_2 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _mstatusNew_WIRE_4_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] _mstatusNew_T_54 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [3:0] next_csr_mstatus_hi_lo_hi_2 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [7:0] next_csr_mstatus_hi_lo_2 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_59 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_WIRE_4_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_58 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_2 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_57 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [2:0] next_csr_mstatus_hi_hi_lo_2 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_62 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [7:0] _mstatusNew_WIRE_4_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [7:0] _mstatusNew_T_61 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_2 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _mstatusNew_WIRE_4_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire  _mstatusNew_T_60 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:55]
  wire [9:0] next_csr_mstatus_hi_hi_hi_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [12:0] next_csr_mstatus_hi_hi_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [20:0] next_csr_mstatus_hi_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [31:0] _next_csr_mstatus_T_2 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _T_622 = 5'h2 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [1:0] _T_623 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:20]
  wire  _T_624 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:27]
  wire [15:0] _next_csr_stval_T = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:69]
  wire [31:0] _next_csr_stval_T_1 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_3181 = inst[1:0] != 2'h3 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:{45,62} 272:41]
  wire  _T_625 = 5'h1 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [1:0] _T_626 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:20]
  wire  _T_627 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:27]
  wire [15:0] _next_csr_stval_T_2 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:69]
  wire [31:0] _next_csr_stval_T_3 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_3182 = _T_624 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 275:{45,62} 276:41]
  wire  _T_628 = 5'h3 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [1:0] _T_629 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:20]
  wire  _T_630 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:27]
  wire [15:0] _next_csr_stval_T_4 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:69]
  wire [31:0] _next_csr_stval_T_5 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_3183 = _T_624 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 280:{45,62} 281:41]
  wire  _T_631 = 5'hb == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire  _T_632 = 5'h6 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire  _T_633 = 5'h4 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire  _T_634 = 5'h0 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] mem_read_addr = io_valid ? _GEN_2422 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_3313 = mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_3184 = 5'h4 == exceptionNO ? mem_read_addr : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 296:26 259:35]
  wire [31:0] mem_write_addr = io_valid ? _GEN_2509 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_3320 = mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_3185 = 5'h6 == exceptionNO ? mem_write_addr : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 292:26]
  wire [31:0] _GEN_3186 = 5'hb == exceptionNO ? 32'h0 : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 288:26]
  wire [31:0] _GEN_3187 = 5'h3 == exceptionNO ? _GEN_3181 : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] _GEN_3188 = 5'h1 == exceptionNO ? _GEN_3181 : _GEN_3187; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] _GEN_3189 = 5'h2 == exceptionNO ? _GEN_3181 : _GEN_3188; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [29:0] _next_pc_T_20 = io_now_csr_stvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:46]
  wire [31:0] _next_pc_T_21 = {io_now_csr_stvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:62]
  wire [29:0] _next_pc_T_22 = io_now_csr_stvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:45]
  wire [31:0] _next_pc_T_23 = {27'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_3345 = {{2'd0}, io_now_csr_stvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [32:0] _next_pc_T_24 = _GEN_3345 + _next_pc_T_23; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [31:0] _next_pc_T_25 = _GEN_3345 + _next_pc_T_23; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [33:0] _next_pc_T_26 = {_next_pc_T_25, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:92]
  wire [33:0] _GEN_3191 = 2'h1 == io_now_csr_stvec[1:0] ? _next_pc_T_26 : {{2'd0}, _GEN_3178}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 317:29]
  wire [33:0] _GEN_3193 = 2'h0 == io_now_csr_stvec[1:0] ? {{2'd0}, _next_pc_T_21} : _GEN_3191; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 312:29]
  wire  _T_638 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] now_csr_scause = io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3194 = 8'h20 == io_now_csr_MXLEN ? _next_csr_scause_T_1 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 252:23]
  wire  _GEN_3199 = 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 165:35 258:35]
  wire [31:0] now_csr_stval = io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3200 = 8'h20 == io_now_csr_MXLEN ? _GEN_3189 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [31:0] _GEN_3201 = 8'h20 == io_now_csr_MXLEN ? _next_csr_mstatus_T_2 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 260:35]
  wire [33:0] _GEN_3203 = 8'h20 == io_now_csr_MXLEN ? _GEN_3193 : {{2'd0}, _GEN_3178}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [30:0] _next_csr_mcause_T = {26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _next_csr_mcause_T_1 = {1'h0,26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 185:41]
  wire [1:0] next_csr_mstatus_lo_lo_lo_3 = {mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_3 = {mstatusOld_pad2,mstatusNew_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [2:0] next_csr_mstatus_lo_lo_hi_3 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [4:0] next_csr_mstatus_lo_lo_3 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_lo_hi_lo_3 = {mstatusOld_ube,mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_3 = {mstatusOld_vs,mstatusNew_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [3:0] next_csr_mstatus_lo_hi_hi_3 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [5:0] next_csr_mstatus_lo_hi_3 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,
    mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [10:0] next_csr_mstatus_lo_3 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,mstatusNew_2_spie
    ,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [3:0] next_csr_mstatus_hi_lo_lo_3 = {mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_3 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [3:0] next_csr_mstatus_hi_lo_hi_3 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [7:0] next_csr_mstatus_hi_lo_3 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_3 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [2:0] next_csr_mstatus_hi_hi_lo_3 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_3 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [9:0] next_csr_mstatus_hi_hi_hi_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [12:0] next_csr_mstatus_hi_hi_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [20:0] next_csr_mstatus_hi_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire [31:0] _next_csr_mstatus_T_3 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 193:38]
  wire  _T_640 = 5'h2 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_641 = 5'h1 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [1:0] _T_642 = inst[1:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:20]
  wire  _T_643 = inst[1:0] != 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:27]
  wire [15:0] _next_csr_mtval_T_18 = inst[15:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:69]
  wire [31:0] _next_csr_mtval_T_19 = inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _GEN_3204 = _T_624 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 204:{45,62} 205:41]
  wire  _T_644 = 5'hb == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_645 = 5'h6 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_646 = 5'h4 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_647 = 5'h0 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_648 = 5'h7 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_649 = 5'hd == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire  _T_650 = 5'hc == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [31:0] _GEN_3205 = _T_633 ? mem_read_addr : 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 192:24 196:29 215:26]
  wire [31:0] _GEN_3206 = _T_632 ? mem_write_addr : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 211:26]
  wire [31:0] _GEN_3207 = _T_631 ? 32'h0 : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 208:26]
  wire [31:0] _GEN_3208 = _T_625 ? _GEN_3181 : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [31:0] _GEN_3209 = _T_622 ? 32'h0 : _GEN_3208; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 199:26]
  wire [29:0] _next_pc_T_27 = io_now_csr_mtvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:46]
  wire [31:0] _next_pc_T_28 = {io_now_csr_mtvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:62]
  wire [29:0] _next_pc_T_29 = io_now_csr_mtvec[31:2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:45]
  wire [31:0] _next_pc_T_30 = {27'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_3346 = {{2'd0}, io_now_csr_mtvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [32:0] _next_pc_T_31 = _GEN_3346 + _next_pc_T_23; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [31:0] _next_pc_T_32 = _GEN_3346 + _next_pc_T_23; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [33:0] _next_pc_T_33 = {_next_pc_T_32, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:92]
  wire [33:0] _GEN_3211 = 2'h1 == io_now_csr_mtvec[1:0] ? _next_pc_T_33 : {{2'd0}, _GEN_3178}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 243:29]
  wire [33:0] _GEN_3213 = 2'h0 == io_now_csr_mtvec[1:0] ? {{2'd0}, _next_pc_T_28} : _GEN_3211; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 238:29]
  wire  _T_654 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] now_csr_mcause = io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3214 = _T_621 ? _next_csr_scause_T_1 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 185:35]
  wire [1:0] _GEN_3219 = 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 175:35 190:35]
  wire [31:0] _GEN_3220 = _T_621 ? _GEN_3209 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_3221 = _T_621 ? _next_csr_mstatus_T_2 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 193:24]
  wire [33:0] _GEN_3223 = _T_621 ? _GEN_3213 : {{2'd0}, _GEN_3178}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [31:0] _GEN_3229 = delegS ? _GEN_3194 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_3246 = raiseExceptionIntr ? _GEN_3229 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_scause = io_valid ? _GEN_3246 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3335 = next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3238 = delegS ? io_now_csr_mcause : _GEN_3214; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_3252 = raiseExceptionIntr ? _GEN_3238 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_mcause = io_valid ? _GEN_3252 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3338 = next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3224 = delegS ? next_csr_scause : next_csr_mcause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 161:35 171:35]
  wire [1:0] _GEN_3228 = delegS ? 2'h1 : 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [31:0] _GEN_3231 = delegS ? _GEN_3200 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [31:0] _GEN_3232 = delegS ? _GEN_3201 : _GEN_3201; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [33:0] _GEN_3234 = delegS ? _GEN_3203 : _GEN_3223; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [31:0] _GEN_3240 = delegS ? _GEN_1925 : _GEN_3220; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [1:0] next_csr_mstatus_lo_lo_lo_4 = {mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_lo_lo_hi_hi_4 = {mstatusOld_pad2,mstatusNew_2_mie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [2:0] next_csr_mstatus_lo_lo_hi_4 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [4:0] next_csr_mstatus_lo_lo_4 = {mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_lo_hi_lo_4 = {mstatusOld_ube,mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [2:0] next_csr_mstatus_lo_hi_hi_hi_4 = {mstatusOld_vs,mstatusNew_2_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [3:0] next_csr_mstatus_lo_hi_hi_4 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [5:0] next_csr_mstatus_lo_hi_4 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,
    mstatusNew_2_spie}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [10:0] next_csr_mstatus_lo_4 = {mstatusOld_vs,mstatusNew_2_spp,mstatusNew_2_mpie,mstatusOld_ube,mstatusNew_2_spie
    ,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [3:0] next_csr_mstatus_hi_lo_lo_4 = {mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_hi_lo_hi_hi_4 = {mstatusOld_sum,mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [3:0] next_csr_mstatus_hi_lo_hi_4 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [7:0] next_csr_mstatus_hi_lo_4 = {mstatusOld_sum,mstatusOld_mprv,mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [1:0] next_csr_mstatus_hi_hi_lo_hi_4 = {mstatusOld_tw,mstatusOld_tvm}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [2:0] next_csr_mstatus_hi_hi_lo_4 = {mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [8:0] next_csr_mstatus_hi_hi_hi_hi_4 = {mstatusOld_sd,mstatusOld_pad0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [9:0] next_csr_mstatus_hi_hi_hi_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [12:0] next_csr_mstatus_hi_hi_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [20:0] next_csr_mstatus_hi_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire [31:0] _next_csr_mstatus_T_4 = {mstatusOld_sd,mstatusOld_pad0,mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,
    mstatusOld_mxr,next_csr_mstatus_hi_lo_2,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 181:36]
  wire  _GEN_3241 = raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [31:0] _event_WIRE_cause = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_3242 = raiseExceptionIntr ? _GEN_3224 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _event_WIRE_exceptionPC = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_3243 = raiseExceptionIntr ? io_now_pc : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 151:25]
  wire [31:0] _event_WIRE_exceptionInst = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_3244 = raiseExceptionIntr ? inst : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 152:25]
  wire [1:0] _GEN_3245 = raiseExceptionIntr ? _GEN_3228 : _GEN_3157; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _GEN_3248 = raiseExceptionIntr ? _GEN_3231 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _GEN_3249 = raiseExceptionIntr ? _next_csr_mstatus_T_2 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 181:22]
  wire [33:0] _GEN_3251 = raiseExceptionIntr ? _GEN_3234 : {{2'd0}, _GEN_3178}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] _GEN_3254 = raiseExceptionIntr ? _GEN_3240 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [31:0] next_csr_cycle = io_valid ? _next_csr_cycle_T_1 : io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 126:20 111:21]
  wire [31:0] _GEN_3258 = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 131:16 115:21]
  wire [2:0] funct3 = io_valid ? _GEN_3174 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 18:24]
  wire [6:0] opcode = io_valid ? _GEN_3176 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 16:24]
  wire [31:0] next_reg_0 = io_valid ? 32'h0 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  wire [31:0] next_reg_1 = io_valid ? _GEN_3087 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_2 = io_valid ? _GEN_3088 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_3 = io_valid ? _GEN_3089 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_4 = io_valid ? _GEN_3090 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_5 = io_valid ? _GEN_3091 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_6 = io_valid ? _GEN_3092 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_7 = io_valid ? _GEN_3093 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_8 = io_valid ? _GEN_3094 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_9 = io_valid ? _GEN_3095 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_10 = io_valid ? _GEN_3096 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_11 = io_valid ? _GEN_3097 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_12 = io_valid ? _GEN_3098 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_13 = io_valid ? _GEN_3099 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_14 = io_valid ? _GEN_3100 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_15 = io_valid ? _GEN_3101 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_16 = io_valid ? _GEN_3102 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_17 = io_valid ? _GEN_3103 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_18 = io_valid ? _GEN_3104 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_19 = io_valid ? _GEN_3105 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_20 = io_valid ? _GEN_3106 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_21 = io_valid ? _GEN_3107 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_22 = io_valid ? _GEN_3108 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_23 = io_valid ? _GEN_3109 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_24 = io_valid ? _GEN_3110 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_25 = io_valid ? _GEN_3111 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_26 = io_valid ? _GEN_3112 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_27 = io_valid ? _GEN_3113 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_28 = io_valid ? _GEN_3114 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_29 = io_valid ? _GEN_3115 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_30 = io_valid ? _GEN_3116 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_reg_31 = io_valid ? _GEN_3117 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [6:0] funct7 = io_valid ? _GEN_3080 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 21:24]
  wire [33:0] _GEN_3305 = io_valid ? _GEN_3251 : {{2'd0}, io_now_pc}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mtval = io_valid ? _GEN_3254 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire  mem_read_valid = io_valid & _GEN_2421; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] mem_read_memWidth = io_valid ? _GEN_2423 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  mem_write_valid = io_valid & _GEN_2508; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] mem_write_memWidth = io_valid ? _GEN_2510 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] mem_write_data = io_valid ? _GEN_2511 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [1:0] next_internal_privilegeMode = io_valid ? _GEN_3245 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mstatus = io_valid ? _GEN_3249 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3330 = retTarget; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _event_WIRE_valid = 1'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire  event_valid = io_valid & raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] event_cause = io_valid ? _GEN_3242 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] event_exceptionPC = io_valid ? _GEN_3243 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] event_exceptionInst = io_valid ? _GEN_3244 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] next_csr_stval = io_valid ? _GEN_3248 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] now_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mstatush = io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mscratch = io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mcounteren = io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mideleg = io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mip = io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_mie = io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_scounteren = io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_sscratch = io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg0 = io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg1 = io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg2 = io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpcfg3 = io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr0 = io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr1 = io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr2 = io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] now_csr_pmpaddr3 = io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] now_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] now_csr_ILEN = io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3265 = next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  wire [31:0] _GEN_3266 = next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3267 = next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3268 = next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3269 = next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3270 = next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3271 = next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3272 = next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3273 = next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3274 = next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3275 = next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3276 = next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3277 = next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3278 = next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3279 = next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3280 = next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3281 = next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3282 = next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3283 = next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3284 = next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3285 = next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3286 = next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3287 = next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3288 = next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3289 = next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3290 = next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3291 = next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3292 = next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3293 = next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3294 = next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3295 = next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3296 = next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_pc = _GEN_3305[31:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 18:18]
  wire [31:0] next_csr_misa = io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3329 = next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_mstatush = io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mscratch = io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mtvec = io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mcounteren = io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mideleg = io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mip = io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_mie = io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3306 = next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] _GEN_3255 = next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 126:20 111:21]
  wire [31:0] next_csr_scounteren = io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] _GEN_3337 = next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] next_csr_sscratch = io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg0 = io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg1 = io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg2 = io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpcfg3 = io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr0 = io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr1 = io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr2 = io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [31:0] next_csr_pmpaddr3 = io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] next_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] next_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [7:0] next_csr_ILEN = io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  wire [1:0] _GEN_3328 = next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [31:0] iFetchpc = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 131:16 115:21]
  wire  _GEN_3312 = mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] _GEN_3314 = mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  _GEN_3319 = mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [5:0] _GEN_3321 = mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [31:0] _GEN_3322 = mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire  _GEN_3331 = event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] _event_WIRE_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] event_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  wire [31:0] _GEN_3332 = event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] _GEN_3333 = event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire [31:0] _GEN_3334 = event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  wire  _exceptionVec_WIRE_10 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  _exceptionVec_WIRE_14 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_10 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire  exceptionVec_14 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:{38,38}]
  wire [6:0] _GEN_3263 = opcode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 16:24]
  wire [2:0] _GEN_3261 = funct3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 18:24]
  wire [6:0] _GEN_3298 = funct7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 21:24]
  wire [1:0] funct2 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 94:{24,24}]
  wire [3:0] funct4 = 4'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 95:{24,24}]
  wire [5:0] funct6 = 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 96:{24,24}]
  wire [1:0] op = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 97:{24,24}]
  wire [2:0] rdP = 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:{24,24}]
  wire [2:0] rs1P = 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:{24,24}]
  wire [2:0] rs2P = 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:{24,24}]
  wire  ph1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:{22,22}]
  wire [4:0] ph5 = 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 103:{52,52}]
  wire [5:0] ph6 = 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 104:{22,22}]
  wire [7:0] ph8 = 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 105:{22,22}]
  wire [2:0] ph3 = 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:{22,22}]
  wire [1:0] ph2 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 106:{52,52}]
  wire [10:0] ph11 = 11'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 107:{22,22}]
  wire [11:0] csrAddr = 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 53:{25,25}]
  wire [31:0] _GEN_3159 = retTarget; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [31:0] _mem_WIRE_read_data = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 119:{22,22}]
  wire  _mstatusOld_WIRE_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [7:0] _mstatusOld_WIRE_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_WIRE_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_20 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [7:0] _mstatusOld_T_19 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_17 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_16 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_15 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_14 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_13 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_12 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_11 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_10 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _mstatusOld_T_9 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_7 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_6 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_4 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_3 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_2 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T_1 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_T = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  _mstatusOld_WIRE_2_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [7:0] _mstatusOld_WIRE_2_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_WIRE_2_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_WIRE_2_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_WIRE_2_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_sie = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_WIRE_2_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_41 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [7:0] _mstatusOld_T_40 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_39 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_38 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_37 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_36 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_35 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_34 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_33 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_32 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusOld_T_30 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_29 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_27 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_26 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_25 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_24 = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_23 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_22 = mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire  _mstatusOld_T_21 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 89:57]
  wire [1:0] _mstatusNew_WIRE_2_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusNew_WIRE_2_mie = mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 90:57]
  wire  _mstatusOld_WIRE_4_sd = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [7:0] _mstatusOld_WIRE_4_pad0 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_tsr = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_tw = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_tvm = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_mxr = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_sum = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_mprv = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_xs = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_fs = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_mpp = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_WIRE_4_vs = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_spp = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_mpie = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_ube = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_spie = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_pad2 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_pad3 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_WIRE_4_pad4 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_62 = mstatusOld_sd; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [7:0] _mstatusOld_T_61 = mstatusOld_pad0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_60 = mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_59 = mstatusOld_tw; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_58 = mstatusOld_tvm; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_57 = mstatusOld_mxr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_56 = mstatusOld_sum; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_55 = mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_54 = mstatusOld_xs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_53 = mstatusOld_fs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_52 = mstatusOld_mpp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire [1:0] _mstatusOld_T_51 = mstatusOld_vs; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_50 = mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_49 = mstatusOld_mpie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_48 = mstatusOld_ube; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_47 = mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_46 = mstatusOld_pad2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_44 = mstatusOld_pad3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  wire  _mstatusOld_T_42 = mstatusOld_pad4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 158:55]
  assign io_iFetchpc = io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 131:16 115:21]
  assign io_mem_read_valid = io_valid & _GEN_2421; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_addr = io_valid ? _GEN_2422 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_memWidth = io_valid ? _GEN_2423 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_valid = io_valid & _GEN_2508; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_addr = io_valid ? _GEN_2509 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_memWidth = io_valid ? _GEN_2510 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_data = io_valid ? _GEN_2511 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_next_reg_0 = io_valid ? 32'h0 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  assign io_next_reg_1 = io_valid ? _GEN_3087 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_2 = io_valid ? _GEN_3088 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_3 = io_valid ? _GEN_3089 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_4 = io_valid ? _GEN_3090 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_5 = io_valid ? _GEN_3091 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_6 = io_valid ? _GEN_3092 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_7 = io_valid ? _GEN_3093 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_8 = io_valid ? _GEN_3094 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_9 = io_valid ? _GEN_3095 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_10 = io_valid ? _GEN_3096 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_11 = io_valid ? _GEN_3097 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_12 = io_valid ? _GEN_3098 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_13 = io_valid ? _GEN_3099 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_14 = io_valid ? _GEN_3100 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_15 = io_valid ? _GEN_3101 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_16 = io_valid ? _GEN_3102 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_17 = io_valid ? _GEN_3103 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_18 = io_valid ? _GEN_3104 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_19 = io_valid ? _GEN_3105 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_20 = io_valid ? _GEN_3106 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_21 = io_valid ? _GEN_3107 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_22 = io_valid ? _GEN_3108 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_23 = io_valid ? _GEN_3109 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_24 = io_valid ? _GEN_3110 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_25 = io_valid ? _GEN_3111 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_26 = io_valid ? _GEN_3112 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_27 = io_valid ? _GEN_3113 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_28 = io_valid ? _GEN_3114 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_29 = io_valid ? _GEN_3115 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_30 = io_valid ? _GEN_3116 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_31 = io_valid ? _GEN_3117 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_pc = _GEN_3305[31:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 18:18]
  assign io_next_csr_misa = io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mstatus = io_valid ? _GEN_3249 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mstatush = io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mscratch = io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mtvec = io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mcounteren = io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mideleg = io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mip = io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mie = io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mepc = io_valid ? _GEN_3253 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mcause = io_valid ? _GEN_3252 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mtval = io_valid ? _GEN_3254 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_cycle = io_valid ? _next_csr_cycle_T_1 : io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 126:20 111:21]
  assign io_next_csr_scounteren = io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_scause = io_valid ? _GEN_3246 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_sepc = io_valid ? _GEN_3247 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_stval = io_valid ? _GEN_3248 : io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_sscratch = io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg0 = io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg1 = io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg2 = io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpcfg3 = io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr0 = io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr1 = io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr2 = io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_pmpaddr3 = io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_ILEN = io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_internal_privilegeMode = io_valid ? _GEN_3245 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_event_valid = io_valid & raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:{36,36}]
  assign io_event_cause = io_valid ? _GEN_3242 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionPC = io_valid ? _GEN_3243 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionInst = io_valid ? _GEN_3244 : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
endmodule
module RiscvCore(
  input         clock,
  input         reset,
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_iFetchpc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_now_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_now_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_now_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_now_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [1:0]  io_now_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mstatush, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mideleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_cycle, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_scounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_stval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_sscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpcfg3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_next_csr_pmpaddr3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_next_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_next_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [7:0]  io_next_csr_ILEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [1:0]  io_next_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [31:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
`endif // RANDOMIZE_REG_INIT
  wire  trans_clock; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_reset; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_iFetchpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [5:0] trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [5:0] trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_intrNO; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [31:0] trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [30:0] _state_state_csr_misaInitVal_T = 31'h40000000; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 335:25]
  wire [8:0] _state_state_csr_misaInitVal_T_1 = 9'h100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire [8:0] _state_state_csr_misaInitVal_T_2 = 9'h100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [12:0] _state_state_csr_misaInitVal_T_3 = 13'h1000; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 320:66]
  wire [12:0] _state_state_csr_misaInitVal_T_4 = 13'h1100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:75]
  wire [30:0] state_state_csr_misaInitVal = 31'h40001100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 341:20]
  wire [31:0] state_state_csr_csr_mstatus = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 353:17]
  wire [31:0] _state_state_csr_mstatusStruct_WIRE = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 353:17]
  wire  _state_state_csr_mstatusStruct_T = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_1 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_2 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_3 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_4 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_5 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_6 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_7 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_8 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_9 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_10 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_11 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] _state_state_csr_mstatusStruct_T_12 = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_13 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_14 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_15 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_16 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_17 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_18 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [7:0] _state_state_csr_mstatusStruct_T_19 = 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  _state_state_csr_mstatusStruct_T_20 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  reg [31:0] state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [31:0] state_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [1:0] state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  wire [31:0] state_state_reg_0 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_1 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_2 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_3 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_4 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_5 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_6 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_7 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_8 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_9 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_10 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_11 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_12 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_13 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_14 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_15 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_16 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_17 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_18 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_19 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_20 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_21 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_22 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_23 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_24 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_25 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_26 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_27 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_28 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_29 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_30 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_reg_31 = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 80:15]
  wire [31:0] state_state_pc = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 78:21 84:15]
  wire [31:0] state_state_csr_csr_misa = 32'h40001100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 343:14]
  wire [31:0] state_state_csr_misa = 32'h40001100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 343:14]
  wire [31:0] state_state_csr_csr_mvendorid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 347:19]
  wire [31:0] state_state_csr_mvendorid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 347:19]
  wire [31:0] state_state_csr_csr_marchid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 349:17]
  wire [31:0] state_state_csr_marchid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 349:17]
  wire [31:0] state_state_csr_csr_mimpid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 351:17]
  wire [31:0] state_state_csr_mimpid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 351:17]
  wire [31:0] state_state_csr_csr_mhartid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 352:17]
  wire [31:0] state_state_csr_mhartid = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 352:17]
  wire [31:0] state_state_csr_mstatus = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 353:17]
  wire [31:0] state_state_csr_csr_mstatush = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 357:20]
  wire [31:0] state_state_csr_mstatush = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 357:20]
  wire [31:0] state_state_csr_csr_mscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 358:20]
  wire [31:0] state_state_csr_mscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 358:20]
  wire [31:0] state_state_csr_csr_mtvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 359:20]
  wire [31:0] state_state_csr_mtvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 359:20]
  wire [31:0] state_state_csr_csr_mcounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 360:20]
  wire [31:0] state_state_csr_mcounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 360:20]
  wire [31:0] state_state_csr_csr_medeleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 361:20]
  wire [31:0] state_state_csr_medeleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 361:20]
  wire [31:0] state_state_csr_csr_mideleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 362:20]
  wire [31:0] state_state_csr_mideleg = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 362:20]
  wire [31:0] state_state_csr_csr_mip = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 363:20]
  wire [31:0] state_state_csr_mip = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 363:20]
  wire [31:0] state_state_csr_csr_mie = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 364:20]
  wire [31:0] state_state_csr_mie = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 364:20]
  wire [31:0] state_state_csr_csr_mepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 365:20]
  wire [31:0] state_state_csr_mepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 365:20]
  wire [31:0] state_state_csr_csr_mcause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 366:20]
  wire [31:0] state_state_csr_mcause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 366:20]
  wire [31:0] state_state_csr_csr_mtval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 367:20]
  wire [31:0] state_state_csr_mtval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 367:20]
  wire [31:0] state_state_csr_csr_cycle = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 368:20]
  wire [31:0] state_state_csr_cycle = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 368:20]
  wire [31:0] state_state_csr_csr_scounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 372:20]
  wire [31:0] state_state_csr_scounteren = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 372:20]
  wire [31:0] state_state_csr_csr_scause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 371:20]
  wire [31:0] state_state_csr_scause = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 371:20]
  wire [31:0] state_state_csr_csr_stvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 373:20]
  wire [31:0] state_state_csr_stvec = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 373:20]
  wire [31:0] state_state_csr_csr_sepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 374:20]
  wire [31:0] state_state_csr_sepc = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 374:20]
  wire [31:0] state_state_csr_csr_stval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 375:20]
  wire [31:0] state_state_csr_stval = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 375:20]
  wire [31:0] state_state_csr_csr_sscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 376:20]
  wire [31:0] state_state_csr_sscratch = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 376:20]
  wire [31:0] state_state_csr_csr_satp = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 378:14]
  wire [31:0] state_state_csr_satp = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 378:14]
  wire [31:0] state_state_csr_csr_pmpcfg0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 386:18]
  wire [31:0] state_state_csr_pmpcfg0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 386:18]
  wire [31:0] state_state_csr_csr_pmpcfg1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 387:18]
  wire [31:0] state_state_csr_pmpcfg1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 387:18]
  wire [31:0] state_state_csr_csr_pmpcfg2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 388:18]
  wire [31:0] state_state_csr_pmpcfg2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 388:18]
  wire [31:0] state_state_csr_csr_pmpcfg3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 389:18]
  wire [31:0] state_state_csr_pmpcfg3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 389:18]
  wire [31:0] state_state_csr_csr_pmpaddr0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 390:18]
  wire [31:0] state_state_csr_pmpaddr0 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 390:18]
  wire [31:0] state_state_csr_csr_pmpaddr1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 391:18]
  wire [31:0] state_state_csr_pmpaddr1 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 391:18]
  wire [31:0] state_state_csr_csr_pmpaddr2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 392:18]
  wire [31:0] state_state_csr_pmpaddr2 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 392:18]
  wire [31:0] state_state_csr_csr_pmpaddr3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 393:18]
  wire [31:0] state_state_csr_pmpaddr3 = 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 393:18]
  wire [7:0] state_state_csr_csr_MXLEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 398:15]
  wire [7:0] state_state_csr_MXLEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 398:15]
  wire [7:0] state_state_csr_csr_IALIGN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 399:16]
  wire [7:0] state_state_csr_IALIGN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 399:16]
  wire [7:0] state_state_csr_csr_ILEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 403:14]
  wire [7:0] state_state_csr_ILEN = 8'h20; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 330:19 403:14]
  wire [1:0] state_state_internal_internal_privilegeMode = 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 61:24 62:28]
  wire [1:0] state_state_internal_privilegeMode = 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 61:24 62:28]
  wire  state_state_csr_mstatusStruct_sd = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [7:0] state_state_csr_mstatusStruct_pad0 = 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_tsr = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_tw = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_tvm = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mxr = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_sum = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mprv = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_xs = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_fs = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_mpp = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire [1:0] state_state_csr_mstatusStruct_vs = 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_spp = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mpie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_ube = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_spie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_pad2 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_mie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_pad3 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_sie = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  wire  state_state_csr_mstatusStruct_pad4 = 1'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 354:45]
  RiscvTrans trans ( // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
    .clock(trans_clock),
    .reset(trans_reset),
    .io_inst(trans_io_inst),
    .io_valid(trans_io_valid),
    .io_iFetchpc(trans_io_iFetchpc),
    .io_mem_read_valid(trans_io_mem_read_valid),
    .io_mem_read_addr(trans_io_mem_read_addr),
    .io_mem_read_memWidth(trans_io_mem_read_memWidth),
    .io_mem_read_data(trans_io_mem_read_data),
    .io_mem_write_valid(trans_io_mem_write_valid),
    .io_mem_write_addr(trans_io_mem_write_addr),
    .io_mem_write_memWidth(trans_io_mem_write_memWidth),
    .io_mem_write_data(trans_io_mem_write_data),
    .io_now_reg_0(trans_io_now_reg_0),
    .io_now_reg_1(trans_io_now_reg_1),
    .io_now_reg_2(trans_io_now_reg_2),
    .io_now_reg_3(trans_io_now_reg_3),
    .io_now_reg_4(trans_io_now_reg_4),
    .io_now_reg_5(trans_io_now_reg_5),
    .io_now_reg_6(trans_io_now_reg_6),
    .io_now_reg_7(trans_io_now_reg_7),
    .io_now_reg_8(trans_io_now_reg_8),
    .io_now_reg_9(trans_io_now_reg_9),
    .io_now_reg_10(trans_io_now_reg_10),
    .io_now_reg_11(trans_io_now_reg_11),
    .io_now_reg_12(trans_io_now_reg_12),
    .io_now_reg_13(trans_io_now_reg_13),
    .io_now_reg_14(trans_io_now_reg_14),
    .io_now_reg_15(trans_io_now_reg_15),
    .io_now_reg_16(trans_io_now_reg_16),
    .io_now_reg_17(trans_io_now_reg_17),
    .io_now_reg_18(trans_io_now_reg_18),
    .io_now_reg_19(trans_io_now_reg_19),
    .io_now_reg_20(trans_io_now_reg_20),
    .io_now_reg_21(trans_io_now_reg_21),
    .io_now_reg_22(trans_io_now_reg_22),
    .io_now_reg_23(trans_io_now_reg_23),
    .io_now_reg_24(trans_io_now_reg_24),
    .io_now_reg_25(trans_io_now_reg_25),
    .io_now_reg_26(trans_io_now_reg_26),
    .io_now_reg_27(trans_io_now_reg_27),
    .io_now_reg_28(trans_io_now_reg_28),
    .io_now_reg_29(trans_io_now_reg_29),
    .io_now_reg_30(trans_io_now_reg_30),
    .io_now_reg_31(trans_io_now_reg_31),
    .io_now_pc(trans_io_now_pc),
    .io_now_csr_misa(trans_io_now_csr_misa),
    .io_now_csr_mvendorid(trans_io_now_csr_mvendorid),
    .io_now_csr_marchid(trans_io_now_csr_marchid),
    .io_now_csr_mimpid(trans_io_now_csr_mimpid),
    .io_now_csr_mhartid(trans_io_now_csr_mhartid),
    .io_now_csr_mstatus(trans_io_now_csr_mstatus),
    .io_now_csr_mstatush(trans_io_now_csr_mstatush),
    .io_now_csr_mscratch(trans_io_now_csr_mscratch),
    .io_now_csr_mtvec(trans_io_now_csr_mtvec),
    .io_now_csr_mcounteren(trans_io_now_csr_mcounteren),
    .io_now_csr_medeleg(trans_io_now_csr_medeleg),
    .io_now_csr_mideleg(trans_io_now_csr_mideleg),
    .io_now_csr_mip(trans_io_now_csr_mip),
    .io_now_csr_mie(trans_io_now_csr_mie),
    .io_now_csr_mepc(trans_io_now_csr_mepc),
    .io_now_csr_mcause(trans_io_now_csr_mcause),
    .io_now_csr_mtval(trans_io_now_csr_mtval),
    .io_now_csr_cycle(trans_io_now_csr_cycle),
    .io_now_csr_scounteren(trans_io_now_csr_scounteren),
    .io_now_csr_scause(trans_io_now_csr_scause),
    .io_now_csr_stvec(trans_io_now_csr_stvec),
    .io_now_csr_sepc(trans_io_now_csr_sepc),
    .io_now_csr_stval(trans_io_now_csr_stval),
    .io_now_csr_sscratch(trans_io_now_csr_sscratch),
    .io_now_csr_satp(trans_io_now_csr_satp),
    .io_now_csr_pmpcfg0(trans_io_now_csr_pmpcfg0),
    .io_now_csr_pmpcfg1(trans_io_now_csr_pmpcfg1),
    .io_now_csr_pmpcfg2(trans_io_now_csr_pmpcfg2),
    .io_now_csr_pmpcfg3(trans_io_now_csr_pmpcfg3),
    .io_now_csr_pmpaddr0(trans_io_now_csr_pmpaddr0),
    .io_now_csr_pmpaddr1(trans_io_now_csr_pmpaddr1),
    .io_now_csr_pmpaddr2(trans_io_now_csr_pmpaddr2),
    .io_now_csr_pmpaddr3(trans_io_now_csr_pmpaddr3),
    .io_now_csr_MXLEN(trans_io_now_csr_MXLEN),
    .io_now_csr_IALIGN(trans_io_now_csr_IALIGN),
    .io_now_csr_ILEN(trans_io_now_csr_ILEN),
    .io_now_internal_privilegeMode(trans_io_now_internal_privilegeMode),
    .io_next_reg_0(trans_io_next_reg_0),
    .io_next_reg_1(trans_io_next_reg_1),
    .io_next_reg_2(trans_io_next_reg_2),
    .io_next_reg_3(trans_io_next_reg_3),
    .io_next_reg_4(trans_io_next_reg_4),
    .io_next_reg_5(trans_io_next_reg_5),
    .io_next_reg_6(trans_io_next_reg_6),
    .io_next_reg_7(trans_io_next_reg_7),
    .io_next_reg_8(trans_io_next_reg_8),
    .io_next_reg_9(trans_io_next_reg_9),
    .io_next_reg_10(trans_io_next_reg_10),
    .io_next_reg_11(trans_io_next_reg_11),
    .io_next_reg_12(trans_io_next_reg_12),
    .io_next_reg_13(trans_io_next_reg_13),
    .io_next_reg_14(trans_io_next_reg_14),
    .io_next_reg_15(trans_io_next_reg_15),
    .io_next_reg_16(trans_io_next_reg_16),
    .io_next_reg_17(trans_io_next_reg_17),
    .io_next_reg_18(trans_io_next_reg_18),
    .io_next_reg_19(trans_io_next_reg_19),
    .io_next_reg_20(trans_io_next_reg_20),
    .io_next_reg_21(trans_io_next_reg_21),
    .io_next_reg_22(trans_io_next_reg_22),
    .io_next_reg_23(trans_io_next_reg_23),
    .io_next_reg_24(trans_io_next_reg_24),
    .io_next_reg_25(trans_io_next_reg_25),
    .io_next_reg_26(trans_io_next_reg_26),
    .io_next_reg_27(trans_io_next_reg_27),
    .io_next_reg_28(trans_io_next_reg_28),
    .io_next_reg_29(trans_io_next_reg_29),
    .io_next_reg_30(trans_io_next_reg_30),
    .io_next_reg_31(trans_io_next_reg_31),
    .io_next_pc(trans_io_next_pc),
    .io_next_csr_misa(trans_io_next_csr_misa),
    .io_next_csr_mvendorid(trans_io_next_csr_mvendorid),
    .io_next_csr_marchid(trans_io_next_csr_marchid),
    .io_next_csr_mimpid(trans_io_next_csr_mimpid),
    .io_next_csr_mhartid(trans_io_next_csr_mhartid),
    .io_next_csr_mstatus(trans_io_next_csr_mstatus),
    .io_next_csr_mstatush(trans_io_next_csr_mstatush),
    .io_next_csr_mscratch(trans_io_next_csr_mscratch),
    .io_next_csr_mtvec(trans_io_next_csr_mtvec),
    .io_next_csr_mcounteren(trans_io_next_csr_mcounteren),
    .io_next_csr_medeleg(trans_io_next_csr_medeleg),
    .io_next_csr_mideleg(trans_io_next_csr_mideleg),
    .io_next_csr_mip(trans_io_next_csr_mip),
    .io_next_csr_mie(trans_io_next_csr_mie),
    .io_next_csr_mepc(trans_io_next_csr_mepc),
    .io_next_csr_mcause(trans_io_next_csr_mcause),
    .io_next_csr_mtval(trans_io_next_csr_mtval),
    .io_next_csr_cycle(trans_io_next_csr_cycle),
    .io_next_csr_scounteren(trans_io_next_csr_scounteren),
    .io_next_csr_scause(trans_io_next_csr_scause),
    .io_next_csr_stvec(trans_io_next_csr_stvec),
    .io_next_csr_sepc(trans_io_next_csr_sepc),
    .io_next_csr_stval(trans_io_next_csr_stval),
    .io_next_csr_sscratch(trans_io_next_csr_sscratch),
    .io_next_csr_satp(trans_io_next_csr_satp),
    .io_next_csr_pmpcfg0(trans_io_next_csr_pmpcfg0),
    .io_next_csr_pmpcfg1(trans_io_next_csr_pmpcfg1),
    .io_next_csr_pmpcfg2(trans_io_next_csr_pmpcfg2),
    .io_next_csr_pmpcfg3(trans_io_next_csr_pmpcfg3),
    .io_next_csr_pmpaddr0(trans_io_next_csr_pmpaddr0),
    .io_next_csr_pmpaddr1(trans_io_next_csr_pmpaddr1),
    .io_next_csr_pmpaddr2(trans_io_next_csr_pmpaddr2),
    .io_next_csr_pmpaddr3(trans_io_next_csr_pmpaddr3),
    .io_next_csr_MXLEN(trans_io_next_csr_MXLEN),
    .io_next_csr_IALIGN(trans_io_next_csr_IALIGN),
    .io_next_csr_ILEN(trans_io_next_csr_ILEN),
    .io_next_internal_privilegeMode(trans_io_next_internal_privilegeMode),
    .io_event_valid(trans_io_event_valid),
    .io_event_intrNO(trans_io_event_intrNO),
    .io_event_cause(trans_io_event_cause),
    .io_event_exceptionPC(trans_io_event_exceptionPC),
    .io_event_exceptionInst(trans_io_event_exceptionInst)
  );
  assign io_iFetchpc = trans_io_iFetchpc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 203:15]
  assign io_mem_read_valid = trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_addr = trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_memWidth = trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_valid = trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_addr = trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_memWidth = trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_data = trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_now_reg_0 = state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_1 = state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_2 = state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_3 = state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_4 = state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_5 = state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_6 = state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_7 = state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_8 = state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_9 = state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_10 = state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_11 = state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_12 = state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_13 = state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_14 = state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_15 = state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_16 = state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_17 = state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_18 = state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_19 = state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_20 = state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_21 = state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_22 = state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_23 = state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_24 = state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_25 = state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_26 = state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_27 = state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_28 = state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_29 = state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_30 = state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_reg_31 = state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_misa = state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mvendorid = state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_marchid = state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mimpid = state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mhartid = state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mstatus = state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mstatush = state_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mscratch = state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mtvec = state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mcounteren = state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_medeleg = state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mideleg = state_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mip = state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mie = state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mepc = state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mcause = state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_mtval = state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_cycle = state_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_scounteren = state_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_scause = state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_stvec = state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_sepc = state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_stval = state_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_sscratch = state_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_satp = state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg0 = state_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg1 = state_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg2 = state_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpcfg3 = state_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr0 = state_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr1 = state_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr2 = state_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_pmpaddr3 = state_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_MXLEN = state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_IALIGN = state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_csr_ILEN = state_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_now_internal_privilegeMode = state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_next_reg_0 = trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_1 = trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_2 = trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_3 = trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_4 = trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_5 = trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_6 = trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_7 = trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_8 = trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_9 = trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_10 = trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_11 = trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_12 = trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_13 = trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_14 = trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_15 = trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_16 = trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_17 = trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_18 = trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_19 = trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_20 = trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_21 = trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_22 = trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_23 = trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_24 = trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_25 = trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_26 = trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_27 = trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_28 = trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_29 = trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_30 = trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_31 = trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_pc = trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_misa = trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mvendorid = trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_marchid = trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mimpid = trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mhartid = trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mstatus = trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mstatush = trans_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mscratch = trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtvec = trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcounteren = trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_medeleg = trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mideleg = trans_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mip = trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mie = trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mepc = trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcause = trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtval = trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_cycle = trans_io_next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_scounteren = trans_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_scause = trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_stvec = trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_sepc = trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_stval = trans_io_next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_sscratch = trans_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_satp = trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg0 = trans_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg1 = trans_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg2 = trans_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpcfg3 = trans_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr0 = trans_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr1 = trans_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr2 = trans_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_pmpaddr3 = trans_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_MXLEN = trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_IALIGN = trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_ILEN = trans_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_internal_privilegeMode = trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_event_valid = trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_intrNO = 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_cause = trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionPC = trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionInst = trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign trans_clock = clock;
  assign trans_reset = reset;
  assign trans_io_inst = io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 192:18]
  assign trans_io_valid = io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 193:18]
  assign trans_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign trans_io_now_reg_0 = state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_1 = state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_2 = state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_3 = state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_4 = state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_5 = state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_6 = state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_7 = state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_8 = state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_9 = state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_10 = state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_11 = state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_12 = state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_13 = state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_14 = state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_15 = state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_16 = state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_17 = state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_18 = state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_19 = state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_20 = state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_21 = state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_22 = state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_23 = state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_24 = state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_25 = state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_26 = state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_27 = state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_28 = state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_29 = state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_30 = state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_31 = state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_misa = state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mvendorid = state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_marchid = state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mimpid = state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mhartid = state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mstatus = state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mstatush = state_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mscratch = state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtvec = state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcounteren = state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_medeleg = state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mideleg = state_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mip = state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mie = state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mepc = state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcause = state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtval = state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_cycle = state_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_scounteren = state_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_scause = state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_stvec = state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_sepc = state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_stval = state_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_sscratch = state_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_satp = state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg0 = state_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg1 = state_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg2 = state_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpcfg3 = state_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr0 = state_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr1 = state_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr2 = state_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_pmpaddr3 = state_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_MXLEN = state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_IALIGN = state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_ILEN = state_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_internal_privilegeMode = state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_0 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_0 <= trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_1 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_1 <= trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_2 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_2 <= trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_3 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_3 <= trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_4 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_4 <= trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_5 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_5 <= trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_6 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_6 <= trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_7 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_7 <= trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_8 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_8 <= trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_9 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_9 <= trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_10 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_10 <= trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_11 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_11 <= trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_12 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_12 <= trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_13 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_13 <= trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_14 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_14 <= trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_15 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_15 <= trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_16 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_16 <= trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_17 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_17 <= trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_18 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_18 <= trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_19 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_19 <= trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_20 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_20 <= trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_21 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_21 <= trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_22 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_22 <= trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_23 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_23 <= trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_24 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_24 <= trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_25 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_25 <= trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_26 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_26 <= trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_27 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_27 <= trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_28 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_28 <= trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_29 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_29 <= trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_30 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_30 <= trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_31 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_31 <= trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_pc <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_pc <= trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_misa <= 32'h40001100; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_misa <= trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mvendorid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mvendorid <= trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_marchid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_marchid <= trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mimpid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mimpid <= trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mhartid <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mhartid <= trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mstatus <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mstatus <= trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mstatush <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mstatush <= trans_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mscratch <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mscratch <= trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtvec <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtvec <= trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcounteren <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcounteren <= trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_medeleg <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_medeleg <= trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mideleg <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mideleg <= trans_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mip <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mip <= trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mie <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mie <= trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mepc <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mepc <= trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcause <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcause <= trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtval <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtval <= trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_cycle <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_cycle <= trans_io_next_csr_cycle; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_scounteren <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_scounteren <= trans_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_scause <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_scause <= trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_stvec <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_stvec <= trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_sepc <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_sepc <= trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_stval <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_stval <= trans_io_next_csr_stval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_sscratch <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_sscratch <= trans_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_satp <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_satp <= trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg0 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg0 <= trans_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg1 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg1 <= trans_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg2 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg2 <= trans_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpcfg3 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpcfg3 <= trans_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr0 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr0 <= trans_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr1 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr1 <= trans_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr2 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr2 <= trans_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_pmpaddr3 <= 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_pmpaddr3 <= trans_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_MXLEN <= 8'h20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_MXLEN <= trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_IALIGN <= 8'h20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_IALIGN <= trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_ILEN <= 8'h20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_ILEN <= trans_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_internal_privilegeMode <= 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_internal_privilegeMode <= trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  state_reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state_reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  state_reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  state_reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  state_reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  state_reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  state_reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  state_reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_reg_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  state_reg_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  state_reg_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  state_reg_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  state_reg_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  state_reg_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  state_reg_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  state_reg_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  state_reg_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  state_reg_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  state_reg_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  state_reg_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  state_reg_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  state_reg_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  state_reg_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  state_reg_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  state_reg_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  state_reg_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  state_reg_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  state_reg_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  state_reg_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  state_reg_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  state_reg_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  state_pc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  state_csr_misa = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  state_csr_mvendorid = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  state_csr_marchid = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  state_csr_mimpid = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  state_csr_mhartid = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  state_csr_mstatus = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  state_csr_mstatush = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  state_csr_mscratch = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  state_csr_mtvec = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  state_csr_mcounteren = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  state_csr_medeleg = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  state_csr_mideleg = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  state_csr_mip = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  state_csr_mie = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  state_csr_mepc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  state_csr_mcause = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  state_csr_mtval = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  state_csr_cycle = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  state_csr_scounteren = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  state_csr_scause = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  state_csr_stvec = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  state_csr_sepc = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  state_csr_stval = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  state_csr_sscratch = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  state_csr_satp = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  state_csr_pmpcfg0 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  state_csr_pmpcfg1 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  state_csr_pmpcfg2 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  state_csr_pmpcfg3 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  state_csr_pmpaddr0 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  state_csr_pmpaddr1 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  state_csr_pmpaddr2 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  state_csr_pmpaddr3 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  state_csr_MXLEN = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  state_csr_IALIGN = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  state_csr_ILEN = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  state_internal_privilegeMode = _RAND_69[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CheckerWithResult(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mstatush, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_medeleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mideleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_cycle, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_scounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_scause, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_stvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_sepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_stval, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_sscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_satp, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg0, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg1, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg2, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpcfg3, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr0, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr1, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr2, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_result_csr_pmpaddr3, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [7:0]  io_result_csr_MXLEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [7:0]  io_result_csr_IALIGN, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [7:0]  io_result_csr_ILEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [1:0]  io_result_internal_privilegeMode, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
  input  [31:0] io_mem_write_data // @[src/main/scala/rvspeccore/checker/Checker.scala 88:16]
);
  wire  specCore_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_iFetchpc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [5:0] specCore_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [5:0] specCore_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_now_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_now_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [1:0] specCore_io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_next_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [7:0] specCore_io_next_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [1:0] specCore_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire [31:0] specCore_io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
  wire  _T = io_mem_read_valid == specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 129:46]
  wire  _T_1 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
  wire  _T_2 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
  wire  _T_3 = ~(io_mem_read_valid == specCore_io_mem_read_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
  wire  _T_4 = io_mem_read_valid | specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 130:43]
  wire  _T_5 = io_mem_read_addr == specCore_io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:47]
  wire  _T_6 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _T_7 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _T_8 = ~(io_mem_read_addr == specCore_io_mem_read_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _T_9 = io_mem_read_memWidth == specCore_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:51]
  wire  _T_10 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _T_11 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _T_12 = ~(io_mem_read_memWidth == specCore_io_mem_read_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _T_13 = io_mem_write_valid == specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 134:47]
  wire  _T_14 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
  wire  _T_15 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
  wire  _T_16 = ~(io_mem_write_valid == specCore_io_mem_write_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
  wire  _T_17 = io_mem_write_valid | specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 135:44]
  wire  _T_18 = io_mem_write_addr == specCore_io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:48]
  wire  _T_19 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _T_20 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _T_21 = ~(io_mem_write_addr == specCore_io_mem_write_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _T_22 = io_mem_write_data == specCore_io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:48]
  wire  _T_23 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _T_24 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _T_25 = ~(io_mem_write_data == specCore_io_mem_write_data); // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _T_26 = io_mem_write_memWidth == specCore_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:52]
  wire  _T_27 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _T_28 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _T_29 = ~(io_mem_write_memWidth == specCore_io_mem_write_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _T_30 = io_instCommit_pc == specCore_io_now_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:39]
  wire  _T_31 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _T_32 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _T_33 = ~(io_instCommit_pc == specCore_io_now_pc); // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _T_34 = io_result_csr_misa == specCore_io_next_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_35 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_36 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_37 = ~(io_result_csr_misa == specCore_io_next_csr_misa); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_38 = io_result_csr_mvendorid == specCore_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_39 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_40 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_41 = ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_42 = io_result_csr_marchid == specCore_io_next_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_43 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_44 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_45 = ~(io_result_csr_marchid == specCore_io_next_csr_marchid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_46 = io_result_csr_mimpid == specCore_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_47 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_48 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_49 = ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_50 = io_result_csr_mhartid == specCore_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_51 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_52 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_53 = ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_54 = io_result_csr_mstatus == specCore_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_55 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_56 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_57 = ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_58 = io_result_csr_mscratch == specCore_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_59 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_60 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_61 = ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_62 = io_result_csr_mtvec == specCore_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_63 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_64 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_65 = ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_66 = io_result_csr_mcounteren == specCore_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_67 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_68 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_69 = ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_70 = io_result_csr_mip == specCore_io_next_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_71 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_72 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_73 = ~(io_result_csr_mip == specCore_io_next_csr_mip); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_74 = io_result_csr_mie == specCore_io_next_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_75 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_76 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_77 = ~(io_result_csr_mie == specCore_io_next_csr_mie); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_78 = io_result_csr_mepc == specCore_io_next_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_79 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_80 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_81 = ~(io_result_csr_mepc == specCore_io_next_csr_mepc); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_82 = io_result_csr_mcause == specCore_io_next_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_83 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_84 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_85 = ~(io_result_csr_mcause == specCore_io_next_csr_mcause); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_86 = io_result_csr_mtval == specCore_io_next_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:40]
  wire  _T_87 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_88 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_89 = ~(io_result_csr_mtval == specCore_io_next_csr_mtval); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _T_90 = io_result_reg_0 == specCore_io_next_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_91 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_92 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_93 = ~(io_result_reg_0 == specCore_io_next_reg_0); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_94 = io_result_reg_1 == specCore_io_next_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_95 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_96 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_97 = ~(io_result_reg_1 == specCore_io_next_reg_1); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_98 = io_result_reg_2 == specCore_io_next_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_99 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_100 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_101 = ~(io_result_reg_2 == specCore_io_next_reg_2); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_102 = io_result_reg_3 == specCore_io_next_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_103 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_104 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_105 = ~(io_result_reg_3 == specCore_io_next_reg_3); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_106 = io_result_reg_4 == specCore_io_next_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_107 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_108 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_109 = ~(io_result_reg_4 == specCore_io_next_reg_4); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_110 = io_result_reg_5 == specCore_io_next_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_111 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_112 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_113 = ~(io_result_reg_5 == specCore_io_next_reg_5); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_114 = io_result_reg_6 == specCore_io_next_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_115 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_116 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_117 = ~(io_result_reg_6 == specCore_io_next_reg_6); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_118 = io_result_reg_7 == specCore_io_next_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_119 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_120 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_121 = ~(io_result_reg_7 == specCore_io_next_reg_7); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_122 = io_result_reg_8 == specCore_io_next_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_123 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_124 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_125 = ~(io_result_reg_8 == specCore_io_next_reg_8); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_126 = io_result_reg_9 == specCore_io_next_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_127 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_128 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_129 = ~(io_result_reg_9 == specCore_io_next_reg_9); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_130 = io_result_reg_10 == specCore_io_next_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_131 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_132 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_133 = ~(io_result_reg_10 == specCore_io_next_reg_10); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_134 = io_result_reg_11 == specCore_io_next_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_135 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_136 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_137 = ~(io_result_reg_11 == specCore_io_next_reg_11); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_138 = io_result_reg_12 == specCore_io_next_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_139 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_140 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_141 = ~(io_result_reg_12 == specCore_io_next_reg_12); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_142 = io_result_reg_13 == specCore_io_next_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_143 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_144 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_145 = ~(io_result_reg_13 == specCore_io_next_reg_13); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_146 = io_result_reg_14 == specCore_io_next_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_147 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_148 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_149 = ~(io_result_reg_14 == specCore_io_next_reg_14); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_150 = io_result_reg_15 == specCore_io_next_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_151 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_152 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_153 = ~(io_result_reg_15 == specCore_io_next_reg_15); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_154 = io_result_reg_16 == specCore_io_next_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_155 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_156 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_157 = ~(io_result_reg_16 == specCore_io_next_reg_16); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_158 = io_result_reg_17 == specCore_io_next_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_159 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_160 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_161 = ~(io_result_reg_17 == specCore_io_next_reg_17); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_162 = io_result_reg_18 == specCore_io_next_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_163 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_164 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_165 = ~(io_result_reg_18 == specCore_io_next_reg_18); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_166 = io_result_reg_19 == specCore_io_next_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_167 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_168 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_169 = ~(io_result_reg_19 == specCore_io_next_reg_19); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_170 = io_result_reg_20 == specCore_io_next_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_171 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_172 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_173 = ~(io_result_reg_20 == specCore_io_next_reg_20); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_174 = io_result_reg_21 == specCore_io_next_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_175 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_176 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_177 = ~(io_result_reg_21 == specCore_io_next_reg_21); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_178 = io_result_reg_22 == specCore_io_next_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_179 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_180 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_181 = ~(io_result_reg_22 == specCore_io_next_reg_22); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_182 = io_result_reg_23 == specCore_io_next_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_183 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_184 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_185 = ~(io_result_reg_23 == specCore_io_next_reg_23); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_186 = io_result_reg_24 == specCore_io_next_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_187 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_188 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_189 = ~(io_result_reg_24 == specCore_io_next_reg_24); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_190 = io_result_reg_25 == specCore_io_next_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_191 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_192 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_193 = ~(io_result_reg_25 == specCore_io_next_reg_25); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_194 = io_result_reg_26 == specCore_io_next_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_195 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_196 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_197 = ~(io_result_reg_26 == specCore_io_next_reg_26); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_198 = io_result_reg_27 == specCore_io_next_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_199 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_200 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_201 = ~(io_result_reg_27 == specCore_io_next_reg_27); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_202 = io_result_reg_28 == specCore_io_next_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_203 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_204 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_205 = ~(io_result_reg_28 == specCore_io_next_reg_28); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_206 = io_result_reg_29 == specCore_io_next_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_207 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_208 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_209 = ~(io_result_reg_29 == specCore_io_next_reg_29); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_210 = io_result_reg_30 == specCore_io_next_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_211 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_212 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_213 = ~(io_result_reg_30 == specCore_io_next_reg_30); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_214 = io_result_reg_31 == specCore_io_next_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:43]
  wire  _T_215 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_216 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_217 = ~(io_result_reg_31 == specCore_io_next_reg_31); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _T_218 = io_event_valid | specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 239:33]
  wire  _T_219 = io_event_valid == specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 241:32]
  wire  _T_220 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _T_221 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _T_222 = ~_T_219; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _T_223 = io_event_intrNO == 32'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:38]
  wire  _T_224 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _T_225 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _T_226 = ~(io_event_intrNO == 32'h0); // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _T_227 = io_event_cause == specCore_io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:37]
  wire  _T_228 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _T_229 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _T_230 = ~(io_event_cause == specCore_io_event_cause); // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _T_231 = io_event_exceptionPC == specCore_io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:43]
  wire  _T_232 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _T_233 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _T_234 = ~(io_event_exceptionPC == specCore_io_event_exceptionPC); // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _T_235 = io_event_exceptionInst == specCore_io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:45]
  wire  _T_236 = reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  wire  _T_237 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  wire  _T_238 = ~(io_event_exceptionInst == specCore_io_event_exceptionInst); // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  wire  _GEN_0 = _T_4 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
  wire  _GEN_1 = _T_4 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
  wire  _GEN_2 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
  wire  _GEN_3 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
  wire  _GEN_4 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
  wire  _GEN_5 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
  wire  _GEN_6 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_7 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_8 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_9 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_10 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_11 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_12 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_13 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_14 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_15 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_16 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_17 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_18 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_19 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
  wire  _GEN_20 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_21 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_22 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_23 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_24 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_25 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_26 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_27 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_28 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_29 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_30 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_31 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_32 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_33 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_34 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_35 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_36 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_37 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_38 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_39 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_40 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_41 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_42 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_43 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_44 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_45 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_46 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_47 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_48 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_49 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_50 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_51 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
  wire  _GEN_52 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
  wire  _GEN_53 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
  wire  _GEN_54 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
  wire  _GEN_55 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
  wire  _GEN_56 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
  RiscvCore specCore ( // @[src/main/scala/rvspeccore/checker/Checker.scala 114:24]
    .clock(specCore_clock),
    .reset(specCore_reset),
    .io_inst(specCore_io_inst),
    .io_valid(specCore_io_valid),
    .io_iFetchpc(specCore_io_iFetchpc),
    .io_mem_read_valid(specCore_io_mem_read_valid),
    .io_mem_read_addr(specCore_io_mem_read_addr),
    .io_mem_read_memWidth(specCore_io_mem_read_memWidth),
    .io_mem_read_data(specCore_io_mem_read_data),
    .io_mem_write_valid(specCore_io_mem_write_valid),
    .io_mem_write_addr(specCore_io_mem_write_addr),
    .io_mem_write_memWidth(specCore_io_mem_write_memWidth),
    .io_mem_write_data(specCore_io_mem_write_data),
    .io_now_reg_0(specCore_io_now_reg_0),
    .io_now_reg_1(specCore_io_now_reg_1),
    .io_now_reg_2(specCore_io_now_reg_2),
    .io_now_reg_3(specCore_io_now_reg_3),
    .io_now_reg_4(specCore_io_now_reg_4),
    .io_now_reg_5(specCore_io_now_reg_5),
    .io_now_reg_6(specCore_io_now_reg_6),
    .io_now_reg_7(specCore_io_now_reg_7),
    .io_now_reg_8(specCore_io_now_reg_8),
    .io_now_reg_9(specCore_io_now_reg_9),
    .io_now_reg_10(specCore_io_now_reg_10),
    .io_now_reg_11(specCore_io_now_reg_11),
    .io_now_reg_12(specCore_io_now_reg_12),
    .io_now_reg_13(specCore_io_now_reg_13),
    .io_now_reg_14(specCore_io_now_reg_14),
    .io_now_reg_15(specCore_io_now_reg_15),
    .io_now_reg_16(specCore_io_now_reg_16),
    .io_now_reg_17(specCore_io_now_reg_17),
    .io_now_reg_18(specCore_io_now_reg_18),
    .io_now_reg_19(specCore_io_now_reg_19),
    .io_now_reg_20(specCore_io_now_reg_20),
    .io_now_reg_21(specCore_io_now_reg_21),
    .io_now_reg_22(specCore_io_now_reg_22),
    .io_now_reg_23(specCore_io_now_reg_23),
    .io_now_reg_24(specCore_io_now_reg_24),
    .io_now_reg_25(specCore_io_now_reg_25),
    .io_now_reg_26(specCore_io_now_reg_26),
    .io_now_reg_27(specCore_io_now_reg_27),
    .io_now_reg_28(specCore_io_now_reg_28),
    .io_now_reg_29(specCore_io_now_reg_29),
    .io_now_reg_30(specCore_io_now_reg_30),
    .io_now_reg_31(specCore_io_now_reg_31),
    .io_now_pc(specCore_io_now_pc),
    .io_now_csr_misa(specCore_io_now_csr_misa),
    .io_now_csr_mvendorid(specCore_io_now_csr_mvendorid),
    .io_now_csr_marchid(specCore_io_now_csr_marchid),
    .io_now_csr_mimpid(specCore_io_now_csr_mimpid),
    .io_now_csr_mhartid(specCore_io_now_csr_mhartid),
    .io_now_csr_mstatus(specCore_io_now_csr_mstatus),
    .io_now_csr_mstatush(specCore_io_now_csr_mstatush),
    .io_now_csr_mscratch(specCore_io_now_csr_mscratch),
    .io_now_csr_mtvec(specCore_io_now_csr_mtvec),
    .io_now_csr_mcounteren(specCore_io_now_csr_mcounteren),
    .io_now_csr_medeleg(specCore_io_now_csr_medeleg),
    .io_now_csr_mideleg(specCore_io_now_csr_mideleg),
    .io_now_csr_mip(specCore_io_now_csr_mip),
    .io_now_csr_mie(specCore_io_now_csr_mie),
    .io_now_csr_mepc(specCore_io_now_csr_mepc),
    .io_now_csr_mcause(specCore_io_now_csr_mcause),
    .io_now_csr_mtval(specCore_io_now_csr_mtval),
    .io_now_csr_cycle(specCore_io_now_csr_cycle),
    .io_now_csr_scounteren(specCore_io_now_csr_scounteren),
    .io_now_csr_scause(specCore_io_now_csr_scause),
    .io_now_csr_stvec(specCore_io_now_csr_stvec),
    .io_now_csr_sepc(specCore_io_now_csr_sepc),
    .io_now_csr_stval(specCore_io_now_csr_stval),
    .io_now_csr_sscratch(specCore_io_now_csr_sscratch),
    .io_now_csr_satp(specCore_io_now_csr_satp),
    .io_now_csr_pmpcfg0(specCore_io_now_csr_pmpcfg0),
    .io_now_csr_pmpcfg1(specCore_io_now_csr_pmpcfg1),
    .io_now_csr_pmpcfg2(specCore_io_now_csr_pmpcfg2),
    .io_now_csr_pmpcfg3(specCore_io_now_csr_pmpcfg3),
    .io_now_csr_pmpaddr0(specCore_io_now_csr_pmpaddr0),
    .io_now_csr_pmpaddr1(specCore_io_now_csr_pmpaddr1),
    .io_now_csr_pmpaddr2(specCore_io_now_csr_pmpaddr2),
    .io_now_csr_pmpaddr3(specCore_io_now_csr_pmpaddr3),
    .io_now_csr_MXLEN(specCore_io_now_csr_MXLEN),
    .io_now_csr_IALIGN(specCore_io_now_csr_IALIGN),
    .io_now_csr_ILEN(specCore_io_now_csr_ILEN),
    .io_now_internal_privilegeMode(specCore_io_now_internal_privilegeMode),
    .io_next_reg_0(specCore_io_next_reg_0),
    .io_next_reg_1(specCore_io_next_reg_1),
    .io_next_reg_2(specCore_io_next_reg_2),
    .io_next_reg_3(specCore_io_next_reg_3),
    .io_next_reg_4(specCore_io_next_reg_4),
    .io_next_reg_5(specCore_io_next_reg_5),
    .io_next_reg_6(specCore_io_next_reg_6),
    .io_next_reg_7(specCore_io_next_reg_7),
    .io_next_reg_8(specCore_io_next_reg_8),
    .io_next_reg_9(specCore_io_next_reg_9),
    .io_next_reg_10(specCore_io_next_reg_10),
    .io_next_reg_11(specCore_io_next_reg_11),
    .io_next_reg_12(specCore_io_next_reg_12),
    .io_next_reg_13(specCore_io_next_reg_13),
    .io_next_reg_14(specCore_io_next_reg_14),
    .io_next_reg_15(specCore_io_next_reg_15),
    .io_next_reg_16(specCore_io_next_reg_16),
    .io_next_reg_17(specCore_io_next_reg_17),
    .io_next_reg_18(specCore_io_next_reg_18),
    .io_next_reg_19(specCore_io_next_reg_19),
    .io_next_reg_20(specCore_io_next_reg_20),
    .io_next_reg_21(specCore_io_next_reg_21),
    .io_next_reg_22(specCore_io_next_reg_22),
    .io_next_reg_23(specCore_io_next_reg_23),
    .io_next_reg_24(specCore_io_next_reg_24),
    .io_next_reg_25(specCore_io_next_reg_25),
    .io_next_reg_26(specCore_io_next_reg_26),
    .io_next_reg_27(specCore_io_next_reg_27),
    .io_next_reg_28(specCore_io_next_reg_28),
    .io_next_reg_29(specCore_io_next_reg_29),
    .io_next_reg_30(specCore_io_next_reg_30),
    .io_next_reg_31(specCore_io_next_reg_31),
    .io_next_pc(specCore_io_next_pc),
    .io_next_csr_misa(specCore_io_next_csr_misa),
    .io_next_csr_mvendorid(specCore_io_next_csr_mvendorid),
    .io_next_csr_marchid(specCore_io_next_csr_marchid),
    .io_next_csr_mimpid(specCore_io_next_csr_mimpid),
    .io_next_csr_mhartid(specCore_io_next_csr_mhartid),
    .io_next_csr_mstatus(specCore_io_next_csr_mstatus),
    .io_next_csr_mstatush(specCore_io_next_csr_mstatush),
    .io_next_csr_mscratch(specCore_io_next_csr_mscratch),
    .io_next_csr_mtvec(specCore_io_next_csr_mtvec),
    .io_next_csr_mcounteren(specCore_io_next_csr_mcounteren),
    .io_next_csr_medeleg(specCore_io_next_csr_medeleg),
    .io_next_csr_mideleg(specCore_io_next_csr_mideleg),
    .io_next_csr_mip(specCore_io_next_csr_mip),
    .io_next_csr_mie(specCore_io_next_csr_mie),
    .io_next_csr_mepc(specCore_io_next_csr_mepc),
    .io_next_csr_mcause(specCore_io_next_csr_mcause),
    .io_next_csr_mtval(specCore_io_next_csr_mtval),
    .io_next_csr_cycle(specCore_io_next_csr_cycle),
    .io_next_csr_scounteren(specCore_io_next_csr_scounteren),
    .io_next_csr_scause(specCore_io_next_csr_scause),
    .io_next_csr_stvec(specCore_io_next_csr_stvec),
    .io_next_csr_sepc(specCore_io_next_csr_sepc),
    .io_next_csr_stval(specCore_io_next_csr_stval),
    .io_next_csr_sscratch(specCore_io_next_csr_sscratch),
    .io_next_csr_satp(specCore_io_next_csr_satp),
    .io_next_csr_pmpcfg0(specCore_io_next_csr_pmpcfg0),
    .io_next_csr_pmpcfg1(specCore_io_next_csr_pmpcfg1),
    .io_next_csr_pmpcfg2(specCore_io_next_csr_pmpcfg2),
    .io_next_csr_pmpcfg3(specCore_io_next_csr_pmpcfg3),
    .io_next_csr_pmpaddr0(specCore_io_next_csr_pmpaddr0),
    .io_next_csr_pmpaddr1(specCore_io_next_csr_pmpaddr1),
    .io_next_csr_pmpaddr2(specCore_io_next_csr_pmpaddr2),
    .io_next_csr_pmpaddr3(specCore_io_next_csr_pmpaddr3),
    .io_next_csr_MXLEN(specCore_io_next_csr_MXLEN),
    .io_next_csr_IALIGN(specCore_io_next_csr_IALIGN),
    .io_next_csr_ILEN(specCore_io_next_csr_ILEN),
    .io_next_internal_privilegeMode(specCore_io_next_internal_privilegeMode),
    .io_event_valid(specCore_io_event_valid),
    .io_event_intrNO(specCore_io_event_intrNO),
    .io_event_cause(specCore_io_event_cause),
    .io_event_exceptionPC(specCore_io_event_exceptionPC),
    .io_event_exceptionInst(specCore_io_event_exceptionInst)
  );
  assign specCore_clock = clock;
  assign specCore_reset = reset;
  assign specCore_io_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 116:21]
  assign specCore_io_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 115:21]
  assign specCore_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 140:33]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_mem_read_valid == specCore_io_mem_read_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:129 assert(regDelay(io.mem.get.read.valid) === regDelay(specCore.io.mem.read.valid))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & _T_2 & ~(io_mem_read_addr == specCore_io_mem_read_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:131 assert(regDelay(io.mem.get.read.addr) === regDelay(specCore.io.mem.read.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_0 & ~(io_mem_read_memWidth == specCore_io_mem_read_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:132 assert(regDelay(io.mem.get.read.memWidth) === regDelay(specCore.io.mem.read.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(io_mem_write_valid == specCore_io_mem_write_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:134 assert(regDelay(io.mem.get.write.valid) === regDelay(specCore.io.mem.write.valid))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17 & _T_2 & ~(io_mem_write_addr == specCore_io_mem_write_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:136 assert(regDelay(io.mem.get.write.addr) === regDelay(specCore.io.mem.write.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2 & ~(io_mem_write_data == specCore_io_mem_write_data)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:137 assert(regDelay(io.mem.get.write.data) === regDelay(specCore.io.mem.write.data))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2 & ~(io_mem_write_memWidth == specCore_io_mem_write_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:138 assert(regDelay(io.mem.get.write.memWidth) === regDelay(specCore.io.mem.write.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_instCommit_valid & _T_2 & ~(io_instCommit_pc == specCore_io_now_pc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:225 assert(regDelay(io.instCommit.pc) === regDelay(specCore.io.now.pc))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_misa == specCore_io_next_csr_misa)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_marchid == specCore_io_next_csr_marchid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mip == specCore_io_next_csr_mip)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mie == specCore_io_next_csr_mie)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mepc == specCore_io_next_csr_mepc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mcause == specCore_io_next_csr_mcause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_csr_mtval == specCore_io_next_csr_mtval)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:230 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_0 == specCore_io_next_reg_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_1 == specCore_io_next_reg_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_2 == specCore_io_next_reg_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_3 == specCore_io_next_reg_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_4 == specCore_io_next_reg_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_5 == specCore_io_next_reg_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_6 == specCore_io_next_reg_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_7 == specCore_io_next_reg_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_8 == specCore_io_next_reg_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_9 == specCore_io_next_reg_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_10 == specCore_io_next_reg_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_11 == specCore_io_next_reg_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_12 == specCore_io_next_reg_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_13 == specCore_io_next_reg_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_14 == specCore_io_next_reg_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_15 == specCore_io_next_reg_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_16 == specCore_io_next_reg_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_17 == specCore_io_next_reg_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_18 == specCore_io_next_reg_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_19 == specCore_io_next_reg_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_20 == specCore_io_next_reg_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_21 == specCore_io_next_reg_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_22 == specCore_io_next_reg_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_23 == specCore_io_next_reg_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_24 == specCore_io_next_reg_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_25 == specCore_io_next_reg_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_26 == specCore_io_next_reg_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_27 == specCore_io_next_reg_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_28 == specCore_io_next_reg_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_29 == specCore_io_next_reg_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_30 == specCore_io_next_reg_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & ~(io_result_reg_31 == specCore_io_next_reg_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:235 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_218 & _T_2 & ~_T_219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Checker.scala:240 assert(\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_intrNO == 32'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:243 assert(regDelay(io.event.intrNO) === regDelay(specCore.io.event.intrNO))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_cause == specCore_io_event_cause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:244 assert(regDelay(io.event.cause) === regDelay(specCore.io.event.cause))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_exceptionPC == specCore_io_event_exceptionPC)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:245 assert(regDelay(io.event.exceptionPC) === regDelay(specCore.io.event.exceptionPC))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & ~(io_event_exceptionInst == specCore_io_event_exceptionInst)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:246 assert(regDelay(io.event.exceptionInst) === regDelay(specCore.io.event.exceptionInst))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(io_mem_read_valid == specCore_io_mem_read_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 129:13]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_mem_read_addr == specCore_io_mem_read_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 131:15]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_mem_read_memWidth == specCore_io_mem_read_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 132:15]
    end
    //
    if (_T_2) begin
      assert(io_mem_write_valid == specCore_io_mem_write_valid); // @[src/main/scala/rvspeccore/checker/Checker.scala 134:13]
    end
    //
    if (_T_17 & _T_2) begin
      assert(io_mem_write_addr == specCore_io_mem_write_addr); // @[src/main/scala/rvspeccore/checker/Checker.scala 136:15]
    end
    //
    if (_T_17 & _T_2) begin
      assert(io_mem_write_data == specCore_io_mem_write_data); // @[src/main/scala/rvspeccore/checker/Checker.scala 137:15]
    end
    //
    if (_T_17 & _T_2) begin
      assert(io_mem_write_memWidth == specCore_io_mem_write_memWidth); // @[src/main/scala/rvspeccore/checker/Checker.scala 138:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_instCommit_pc == io_instCommit_pc); // @[src/main/scala/rvspeccore/checker/Checker.scala 225:11]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_misa == specCore_io_next_csr_misa); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_marchid == specCore_io_next_csr_marchid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mimpid == specCore_io_next_csr_mimpid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mhartid == specCore_io_next_csr_mhartid); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mstatus == specCore_io_next_csr_mstatus); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mscratch == specCore_io_next_csr_mscratch); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mtvec == specCore_io_next_csr_mtvec); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mip == specCore_io_next_csr_mip); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mie == specCore_io_next_csr_mie); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mepc == specCore_io_next_csr_mepc); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mcause == specCore_io_next_csr_mcause); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_csr_mtval == specCore_io_next_csr_mtval); // @[src/main/scala/rvspeccore/checker/Checker.scala 230:15]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_0 == specCore_io_next_reg_0); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_1 == io_result_reg_1); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_2 == specCore_io_next_reg_2); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_3 == specCore_io_next_reg_3); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_4 == specCore_io_next_reg_4); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_5 == specCore_io_next_reg_5); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_6 == specCore_io_next_reg_6); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_7 == specCore_io_next_reg_7); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_8 == specCore_io_next_reg_8); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_9 == specCore_io_next_reg_9); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_10 == specCore_io_next_reg_10); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_11 == specCore_io_next_reg_11); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_12 == specCore_io_next_reg_12); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_13 == specCore_io_next_reg_13); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_14 == specCore_io_next_reg_14); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_15 == specCore_io_next_reg_15); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_16 == specCore_io_next_reg_16); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_17 == specCore_io_next_reg_17); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_18 == specCore_io_next_reg_18); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_19 == specCore_io_next_reg_19); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_20 == specCore_io_next_reg_20); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_21 == specCore_io_next_reg_21); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_22 == specCore_io_next_reg_22); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_23 == specCore_io_next_reg_23); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_24 == specCore_io_next_reg_24); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_25 == specCore_io_next_reg_25); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_26 == specCore_io_next_reg_26); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_27 == specCore_io_next_reg_27); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_28 == specCore_io_next_reg_28); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_29 == specCore_io_next_reg_29); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_30 == specCore_io_next_reg_30); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (io_instCommit_valid & _T_2) begin
      assert(io_result_reg_31 == specCore_io_next_reg_31); // @[src/main/scala/rvspeccore/checker/Checker.scala 235:13]
    end
    //
    if (_T_218 & _T_2) begin
      assert(_T_219); // @[src/main/scala/rvspeccore/checker/Checker.scala 240:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_intrNO == 32'h0); // @[src/main/scala/rvspeccore/checker/Checker.scala 243:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_cause == specCore_io_event_cause); // @[src/main/scala/rvspeccore/checker/Checker.scala 244:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_exceptionPC == specCore_io_event_exceptionPC); // @[src/main/scala/rvspeccore/checker/Checker.scala 245:11]
    end
    //
    if (_T_218 & _T_2) begin
      assert(io_event_exceptionInst == specCore_io_event_exceptionInst); // @[src/main/scala/rvspeccore/checker/Checker.scala 246:11]
    end
  end
endmodule
module CheckerWrapper(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mstatush, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_medeleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mideleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_cycle, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_scounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_scause, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_stvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_sepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_stval, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_sscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_satp, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg0, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg1, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg2, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpcfg3, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr0, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr1, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr2, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_result_csr_pmpaddr3, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [7:0]  io_result_csr_MXLEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [7:0]  io_result_csr_IALIGN, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [7:0]  io_result_csr_ILEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [1:0]  io_result_internal_privilegeMode, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [5:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [5:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
  input  [31:0] io_mem_write_data // @[src/main/scala/rvspeccore/checker/Checker.scala 345:14]
);
  wire  checker__clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_instCommit_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_result_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [7:0] checker__io_result_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [7:0] checker__io_result_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [7:0] checker__io_result_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [1:0] checker__io_result_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [5:0] checker__io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire  checker__io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [5:0] checker__io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  wire [31:0] checker__io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
  CheckerWithResult checker_ ( // @[src/main/scala/rvspeccore/checker/Checker.scala 358:23]
    .clock(checker__clock),
    .reset(checker__reset),
    .io_instCommit_valid(checker__io_instCommit_valid),
    .io_instCommit_inst(checker__io_instCommit_inst),
    .io_instCommit_pc(checker__io_instCommit_pc),
    .io_result_reg_0(checker__io_result_reg_0),
    .io_result_reg_1(checker__io_result_reg_1),
    .io_result_reg_2(checker__io_result_reg_2),
    .io_result_reg_3(checker__io_result_reg_3),
    .io_result_reg_4(checker__io_result_reg_4),
    .io_result_reg_5(checker__io_result_reg_5),
    .io_result_reg_6(checker__io_result_reg_6),
    .io_result_reg_7(checker__io_result_reg_7),
    .io_result_reg_8(checker__io_result_reg_8),
    .io_result_reg_9(checker__io_result_reg_9),
    .io_result_reg_10(checker__io_result_reg_10),
    .io_result_reg_11(checker__io_result_reg_11),
    .io_result_reg_12(checker__io_result_reg_12),
    .io_result_reg_13(checker__io_result_reg_13),
    .io_result_reg_14(checker__io_result_reg_14),
    .io_result_reg_15(checker__io_result_reg_15),
    .io_result_reg_16(checker__io_result_reg_16),
    .io_result_reg_17(checker__io_result_reg_17),
    .io_result_reg_18(checker__io_result_reg_18),
    .io_result_reg_19(checker__io_result_reg_19),
    .io_result_reg_20(checker__io_result_reg_20),
    .io_result_reg_21(checker__io_result_reg_21),
    .io_result_reg_22(checker__io_result_reg_22),
    .io_result_reg_23(checker__io_result_reg_23),
    .io_result_reg_24(checker__io_result_reg_24),
    .io_result_reg_25(checker__io_result_reg_25),
    .io_result_reg_26(checker__io_result_reg_26),
    .io_result_reg_27(checker__io_result_reg_27),
    .io_result_reg_28(checker__io_result_reg_28),
    .io_result_reg_29(checker__io_result_reg_29),
    .io_result_reg_30(checker__io_result_reg_30),
    .io_result_reg_31(checker__io_result_reg_31),
    .io_result_pc(checker__io_result_pc),
    .io_result_csr_misa(checker__io_result_csr_misa),
    .io_result_csr_mvendorid(checker__io_result_csr_mvendorid),
    .io_result_csr_marchid(checker__io_result_csr_marchid),
    .io_result_csr_mimpid(checker__io_result_csr_mimpid),
    .io_result_csr_mhartid(checker__io_result_csr_mhartid),
    .io_result_csr_mstatus(checker__io_result_csr_mstatus),
    .io_result_csr_mstatush(checker__io_result_csr_mstatush),
    .io_result_csr_mscratch(checker__io_result_csr_mscratch),
    .io_result_csr_mtvec(checker__io_result_csr_mtvec),
    .io_result_csr_mcounteren(checker__io_result_csr_mcounteren),
    .io_result_csr_medeleg(checker__io_result_csr_medeleg),
    .io_result_csr_mideleg(checker__io_result_csr_mideleg),
    .io_result_csr_mip(checker__io_result_csr_mip),
    .io_result_csr_mie(checker__io_result_csr_mie),
    .io_result_csr_mepc(checker__io_result_csr_mepc),
    .io_result_csr_mcause(checker__io_result_csr_mcause),
    .io_result_csr_mtval(checker__io_result_csr_mtval),
    .io_result_csr_cycle(checker__io_result_csr_cycle),
    .io_result_csr_scounteren(checker__io_result_csr_scounteren),
    .io_result_csr_scause(checker__io_result_csr_scause),
    .io_result_csr_stvec(checker__io_result_csr_stvec),
    .io_result_csr_sepc(checker__io_result_csr_sepc),
    .io_result_csr_stval(checker__io_result_csr_stval),
    .io_result_csr_sscratch(checker__io_result_csr_sscratch),
    .io_result_csr_satp(checker__io_result_csr_satp),
    .io_result_csr_pmpcfg0(checker__io_result_csr_pmpcfg0),
    .io_result_csr_pmpcfg1(checker__io_result_csr_pmpcfg1),
    .io_result_csr_pmpcfg2(checker__io_result_csr_pmpcfg2),
    .io_result_csr_pmpcfg3(checker__io_result_csr_pmpcfg3),
    .io_result_csr_pmpaddr0(checker__io_result_csr_pmpaddr0),
    .io_result_csr_pmpaddr1(checker__io_result_csr_pmpaddr1),
    .io_result_csr_pmpaddr2(checker__io_result_csr_pmpaddr2),
    .io_result_csr_pmpaddr3(checker__io_result_csr_pmpaddr3),
    .io_result_csr_MXLEN(checker__io_result_csr_MXLEN),
    .io_result_csr_IALIGN(checker__io_result_csr_IALIGN),
    .io_result_csr_ILEN(checker__io_result_csr_ILEN),
    .io_result_internal_privilegeMode(checker__io_result_internal_privilegeMode),
    .io_event_valid(checker__io_event_valid),
    .io_event_intrNO(checker__io_event_intrNO),
    .io_event_cause(checker__io_event_cause),
    .io_event_exceptionPC(checker__io_event_exceptionPC),
    .io_event_exceptionInst(checker__io_event_exceptionInst),
    .io_mem_read_valid(checker__io_mem_read_valid),
    .io_mem_read_addr(checker__io_mem_read_addr),
    .io_mem_read_memWidth(checker__io_mem_read_memWidth),
    .io_mem_read_data(checker__io_mem_read_data),
    .io_mem_write_valid(checker__io_mem_write_valid),
    .io_mem_write_addr(checker__io_mem_write_addr),
    .io_mem_write_memWidth(checker__io_mem_write_memWidth),
    .io_mem_write_data(checker__io_mem_write_data)
  );
  assign checker__clock = clock;
  assign checker__reset = reset;
  assign checker__io_instCommit_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 361:25]
  assign checker__io_instCommit_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 361:25]
  assign checker__io_instCommit_pc = io_instCommit_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 361:25]
  assign checker__io_result_reg_0 = io_result_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_1 = io_result_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_2 = io_result_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_3 = io_result_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_4 = io_result_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_5 = io_result_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_6 = io_result_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_7 = io_result_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_8 = io_result_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_9 = io_result_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_10 = io_result_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_11 = io_result_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_12 = io_result_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_13 = io_result_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_14 = io_result_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_15 = io_result_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_16 = io_result_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_17 = io_result_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_18 = io_result_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_19 = io_result_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_20 = io_result_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_21 = io_result_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_22 = io_result_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_23 = io_result_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_24 = io_result_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_25 = io_result_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_26 = io_result_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_27 = io_result_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_28 = io_result_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_29 = io_result_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_30 = io_result_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_reg_31 = io_result_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_pc = io_result_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_misa = io_result_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mvendorid = io_result_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_marchid = io_result_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mimpid = io_result_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mhartid = io_result_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mstatus = io_result_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mstatush = io_result_csr_mstatush; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mscratch = io_result_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mtvec = io_result_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mcounteren = io_result_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_medeleg = io_result_csr_medeleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mideleg = io_result_csr_mideleg; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mip = io_result_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mie = io_result_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mepc = io_result_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mcause = io_result_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_mtval = io_result_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_cycle = io_result_csr_cycle; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_scounteren = io_result_csr_scounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_scause = io_result_csr_scause; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_stvec = io_result_csr_stvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_sepc = io_result_csr_sepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_stval = io_result_csr_stval; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_sscratch = io_result_csr_sscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_satp = io_result_csr_satp; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg0 = io_result_csr_pmpcfg0; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg1 = io_result_csr_pmpcfg1; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg2 = io_result_csr_pmpcfg2; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpcfg3 = io_result_csr_pmpcfg3; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr0 = io_result_csr_pmpaddr0; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr1 = io_result_csr_pmpaddr1; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr2 = io_result_csr_pmpaddr2; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_pmpaddr3 = io_result_csr_pmpaddr3; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_MXLEN = io_result_csr_MXLEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_IALIGN = io_result_csr_IALIGN; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_csr_ILEN = io_result_csr_ILEN; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_result_internal_privilegeMode = io_result_internal_privilegeMode; // @[src/main/scala/rvspeccore/checker/Checker.scala 362:25]
  assign checker__io_event_valid = io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_intrNO = io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_cause = io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_exceptionPC = io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_event_exceptionInst = io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 363:25]
  assign checker__io_mem_read_valid = io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_read_addr = io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_read_memWidth = io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_valid = io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_addr = io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_memWidth = io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
  assign checker__io_mem_write_data = io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 366:24]
endmodule
